magic
tech sky130A
timestamp 1654898173
<< checkpaint >>
rect 9253 12469 11077 14238
rect 570 6652 2479 8638
rect 1661 4930 3123 6476
rect -630 -630 631 631
<< nwell >>
rect -719 14513 10281 17957
rect -719 14457 10285 14513
rect 9737 14013 10285 14457
rect 9863 12753 10317 12754
rect 9781 12262 10317 12753
rect -683 8762 10317 12262
<< nmos >>
rect 49 5851 149 7044
rect 449 5851 549 7044
rect 849 5851 949 7044
rect 1249 5851 1349 7044
rect 1649 5851 1749 7044
<< pmos >>
rect -11 14707 89 17707
rect 489 14707 589 17707
rect 989 14707 1089 17707
rect 1489 14707 1589 17707
rect 1989 14707 2089 17707
rect 2489 14707 2589 17707
rect 2989 14707 3089 17707
rect 3489 14707 3589 17707
rect 3989 14707 4089 17707
rect 4489 14707 4589 17707
rect 4989 14707 5089 17707
rect 5489 14707 5589 17707
rect 5989 14707 6089 17707
rect 6489 14707 6589 17707
rect 6989 14707 7089 17707
rect 7489 14707 7589 17707
rect 7989 14707 8089 17707
rect 8489 14707 8589 17707
rect 8989 14707 9089 17707
rect 9489 14707 9589 17707
rect 9 9012 109 12012
rect 509 9012 609 12012
rect 1009 9012 1109 12012
rect 1509 9012 1609 12012
rect 2009 9012 2109 12012
rect 2509 9012 2609 12012
rect 3009 9012 3109 12012
rect 3509 9012 3609 12012
rect 4009 9012 4109 12012
rect 4509 9012 4609 12012
rect 5009 9012 5109 12012
rect 5509 9012 5609 12012
rect 6009 9012 6109 12012
rect 6509 9012 6609 12012
rect 7009 9012 7109 12012
rect 7509 9012 7609 12012
rect 8009 9012 8109 12012
rect 8509 9012 8609 12012
rect 9009 9012 9109 12012
rect 9509 9012 9609 12012
<< ndiff >>
rect -146 6857 49 7044
rect -146 6757 -104 6857
rect 16 6757 49 6857
rect -146 6657 49 6757
rect -146 6557 -104 6657
rect 16 6557 49 6657
rect -146 6457 49 6557
rect -146 6357 -104 6457
rect 16 6357 49 6457
rect -146 6257 49 6357
rect -146 6157 -104 6257
rect 16 6157 49 6257
rect -146 6057 49 6157
rect -146 5957 -104 6057
rect 16 5957 49 6057
rect -146 5851 49 5957
rect 149 6857 449 7044
rect 149 6757 242 6857
rect 362 6757 449 6857
rect 149 6657 449 6757
rect 149 6557 242 6657
rect 362 6557 449 6657
rect 149 6457 449 6557
rect 149 6357 242 6457
rect 362 6357 449 6457
rect 149 6257 449 6357
rect 149 6157 242 6257
rect 362 6157 449 6257
rect 149 6057 449 6157
rect 149 5957 242 6057
rect 362 5957 449 6057
rect 149 5851 449 5957
rect 549 6857 849 7044
rect 549 6757 648 6857
rect 768 6757 849 6857
rect 549 6657 849 6757
rect 549 6557 648 6657
rect 768 6557 849 6657
rect 549 6457 849 6557
rect 549 6357 648 6457
rect 768 6357 849 6457
rect 549 6257 849 6357
rect 549 6157 648 6257
rect 768 6157 849 6257
rect 549 6057 849 6157
rect 549 5957 648 6057
rect 768 5957 849 6057
rect 549 5851 849 5957
rect 949 6857 1249 7044
rect 949 6757 1018 6857
rect 1138 6757 1249 6857
rect 949 6657 1249 6757
rect 949 6557 1018 6657
rect 1138 6557 1249 6657
rect 949 6457 1249 6557
rect 949 6357 1018 6457
rect 1138 6357 1249 6457
rect 949 6257 1249 6357
rect 949 6157 1018 6257
rect 1138 6157 1249 6257
rect 949 6057 1249 6157
rect 949 5957 1018 6057
rect 1138 5957 1249 6057
rect 949 5851 1249 5957
rect 1349 6857 1649 7044
rect 1349 6757 1424 6857
rect 1544 6757 1649 6857
rect 1349 6657 1649 6757
rect 1349 6557 1424 6657
rect 1544 6557 1649 6657
rect 1349 6457 1649 6557
rect 1349 6357 1424 6457
rect 1544 6357 1649 6457
rect 1349 6257 1649 6357
rect 1349 6157 1424 6257
rect 1544 6157 1649 6257
rect 1349 6057 1649 6157
rect 1349 5957 1424 6057
rect 1544 5957 1649 6057
rect 1349 5851 1649 5957
rect 1749 6857 1905 7044
rect 1749 6757 1770 6857
rect 1890 6757 1905 6857
rect 1749 6657 1905 6757
rect 1749 6557 1770 6657
rect 1890 6557 1905 6657
rect 1749 6457 1905 6557
rect 1749 6357 1770 6457
rect 1890 6357 1905 6457
rect 1749 6257 1905 6357
rect 1749 6157 1770 6257
rect 1890 6157 1905 6257
rect 1749 6057 1905 6157
rect 1749 5957 1770 6057
rect 1890 5957 1905 6057
rect 1749 5851 1905 5957
<< pdiff >>
rect -469 17477 -11 17707
rect -469 17377 -284 17477
rect -184 17377 -11 17477
rect -469 17277 -11 17377
rect -469 17177 -284 17277
rect -184 17177 -11 17277
rect -469 17077 -11 17177
rect -469 16977 -284 17077
rect -184 16977 -11 17077
rect -469 16877 -11 16977
rect -469 16777 -284 16877
rect -184 16777 -11 16877
rect -469 16677 -11 16777
rect -469 16577 -284 16677
rect -184 16577 -11 16677
rect -469 16477 -11 16577
rect -469 16377 -284 16477
rect -184 16377 -11 16477
rect -469 16277 -11 16377
rect -469 16177 -284 16277
rect -184 16177 -11 16277
rect -469 16077 -11 16177
rect -469 15977 -284 16077
rect -184 15977 -11 16077
rect -469 15877 -11 15977
rect -469 15777 -284 15877
rect -184 15777 -11 15877
rect -469 15677 -11 15777
rect -469 15577 -284 15677
rect -184 15577 -11 15677
rect -469 15477 -11 15577
rect -469 15377 -284 15477
rect -184 15377 -11 15477
rect -469 15277 -11 15377
rect -469 15177 -284 15277
rect -184 15177 -11 15277
rect -469 15077 -11 15177
rect -469 14977 -284 15077
rect -184 14977 -11 15077
rect -469 14707 -11 14977
rect 89 17473 489 17707
rect 89 17373 235 17473
rect 335 17373 489 17473
rect 89 17273 489 17373
rect 89 17173 235 17273
rect 335 17173 489 17273
rect 89 17073 489 17173
rect 89 16973 235 17073
rect 335 16973 489 17073
rect 89 16873 489 16973
rect 89 16773 235 16873
rect 335 16773 489 16873
rect 89 16673 489 16773
rect 89 16573 235 16673
rect 335 16573 489 16673
rect 89 16473 489 16573
rect 89 16373 235 16473
rect 335 16373 489 16473
rect 89 16273 489 16373
rect 89 16173 235 16273
rect 335 16173 489 16273
rect 89 16073 489 16173
rect 89 15973 235 16073
rect 335 15973 489 16073
rect 89 15873 489 15973
rect 89 15773 235 15873
rect 335 15773 489 15873
rect 89 15673 489 15773
rect 89 15573 235 15673
rect 335 15573 489 15673
rect 89 15473 489 15573
rect 89 15373 235 15473
rect 335 15373 489 15473
rect 89 15273 489 15373
rect 89 15173 235 15273
rect 335 15173 489 15273
rect 89 15073 489 15173
rect 89 14973 235 15073
rect 335 14973 489 15073
rect 89 14707 489 14973
rect 589 17473 989 17707
rect 589 17373 740 17473
rect 840 17373 989 17473
rect 589 17273 989 17373
rect 589 17173 740 17273
rect 840 17173 989 17273
rect 589 17073 989 17173
rect 589 16973 740 17073
rect 840 16973 989 17073
rect 589 16873 989 16973
rect 589 16773 740 16873
rect 840 16773 989 16873
rect 589 16673 989 16773
rect 589 16573 740 16673
rect 840 16573 989 16673
rect 589 16473 989 16573
rect 589 16373 740 16473
rect 840 16373 989 16473
rect 589 16273 989 16373
rect 589 16173 740 16273
rect 840 16173 989 16273
rect 589 16073 989 16173
rect 589 15973 740 16073
rect 840 15973 989 16073
rect 589 15873 989 15973
rect 589 15773 740 15873
rect 840 15773 989 15873
rect 589 15673 989 15773
rect 589 15573 740 15673
rect 840 15573 989 15673
rect 589 15473 989 15573
rect 589 15373 740 15473
rect 840 15373 989 15473
rect 589 15273 989 15373
rect 589 15173 740 15273
rect 840 15173 989 15273
rect 589 15073 989 15173
rect 589 14973 740 15073
rect 840 14973 989 15073
rect 589 14707 989 14973
rect 1089 17473 1489 17707
rect 1089 17373 1235 17473
rect 1335 17373 1489 17473
rect 1089 17273 1489 17373
rect 1089 17173 1235 17273
rect 1335 17173 1489 17273
rect 1089 17073 1489 17173
rect 1089 16973 1235 17073
rect 1335 16973 1489 17073
rect 1089 16873 1489 16973
rect 1089 16773 1235 16873
rect 1335 16773 1489 16873
rect 1089 16673 1489 16773
rect 1089 16573 1235 16673
rect 1335 16573 1489 16673
rect 1089 16473 1489 16573
rect 1089 16373 1235 16473
rect 1335 16373 1489 16473
rect 1089 16273 1489 16373
rect 1089 16173 1235 16273
rect 1335 16173 1489 16273
rect 1089 16073 1489 16173
rect 1089 15973 1235 16073
rect 1335 15973 1489 16073
rect 1089 15873 1489 15973
rect 1089 15773 1235 15873
rect 1335 15773 1489 15873
rect 1089 15673 1489 15773
rect 1089 15573 1235 15673
rect 1335 15573 1489 15673
rect 1089 15473 1489 15573
rect 1089 15373 1235 15473
rect 1335 15373 1489 15473
rect 1089 15273 1489 15373
rect 1089 15173 1235 15273
rect 1335 15173 1489 15273
rect 1089 15073 1489 15173
rect 1089 14973 1235 15073
rect 1335 14973 1489 15073
rect 1089 14707 1489 14973
rect 1589 17473 1989 17707
rect 1589 17373 1740 17473
rect 1840 17373 1989 17473
rect 1589 17273 1989 17373
rect 1589 17173 1740 17273
rect 1840 17173 1989 17273
rect 1589 17073 1989 17173
rect 1589 16973 1740 17073
rect 1840 16973 1989 17073
rect 1589 16873 1989 16973
rect 1589 16773 1740 16873
rect 1840 16773 1989 16873
rect 1589 16673 1989 16773
rect 1589 16573 1740 16673
rect 1840 16573 1989 16673
rect 1589 16473 1989 16573
rect 1589 16373 1740 16473
rect 1840 16373 1989 16473
rect 1589 16273 1989 16373
rect 1589 16173 1740 16273
rect 1840 16173 1989 16273
rect 1589 16073 1989 16173
rect 1589 15973 1740 16073
rect 1840 15973 1989 16073
rect 1589 15873 1989 15973
rect 1589 15773 1740 15873
rect 1840 15773 1989 15873
rect 1589 15673 1989 15773
rect 1589 15573 1740 15673
rect 1840 15573 1989 15673
rect 1589 15473 1989 15573
rect 1589 15373 1740 15473
rect 1840 15373 1989 15473
rect 1589 15273 1989 15373
rect 1589 15173 1740 15273
rect 1840 15173 1989 15273
rect 1589 15073 1989 15173
rect 1589 14973 1740 15073
rect 1840 14973 1989 15073
rect 1589 14707 1989 14973
rect 2089 17473 2489 17707
rect 2089 17373 2235 17473
rect 2335 17373 2489 17473
rect 2089 17273 2489 17373
rect 2089 17173 2235 17273
rect 2335 17173 2489 17273
rect 2089 17073 2489 17173
rect 2089 16973 2235 17073
rect 2335 16973 2489 17073
rect 2089 16873 2489 16973
rect 2089 16773 2235 16873
rect 2335 16773 2489 16873
rect 2089 16673 2489 16773
rect 2089 16573 2235 16673
rect 2335 16573 2489 16673
rect 2089 16473 2489 16573
rect 2089 16373 2235 16473
rect 2335 16373 2489 16473
rect 2089 16273 2489 16373
rect 2089 16173 2235 16273
rect 2335 16173 2489 16273
rect 2089 16073 2489 16173
rect 2089 15973 2235 16073
rect 2335 15973 2489 16073
rect 2089 15873 2489 15973
rect 2089 15773 2235 15873
rect 2335 15773 2489 15873
rect 2089 15673 2489 15773
rect 2089 15573 2235 15673
rect 2335 15573 2489 15673
rect 2089 15473 2489 15573
rect 2089 15373 2235 15473
rect 2335 15373 2489 15473
rect 2089 15273 2489 15373
rect 2089 15173 2235 15273
rect 2335 15173 2489 15273
rect 2089 15073 2489 15173
rect 2089 14973 2235 15073
rect 2335 14973 2489 15073
rect 2089 14707 2489 14973
rect 2589 17473 2989 17707
rect 2589 17373 2740 17473
rect 2840 17373 2989 17473
rect 2589 17273 2989 17373
rect 2589 17173 2740 17273
rect 2840 17173 2989 17273
rect 2589 17073 2989 17173
rect 2589 16973 2740 17073
rect 2840 16973 2989 17073
rect 2589 16873 2989 16973
rect 2589 16773 2740 16873
rect 2840 16773 2989 16873
rect 2589 16673 2989 16773
rect 2589 16573 2740 16673
rect 2840 16573 2989 16673
rect 2589 16473 2989 16573
rect 2589 16373 2740 16473
rect 2840 16373 2989 16473
rect 2589 16273 2989 16373
rect 2589 16173 2740 16273
rect 2840 16173 2989 16273
rect 2589 16073 2989 16173
rect 2589 15973 2740 16073
rect 2840 15973 2989 16073
rect 2589 15873 2989 15973
rect 2589 15773 2740 15873
rect 2840 15773 2989 15873
rect 2589 15673 2989 15773
rect 2589 15573 2740 15673
rect 2840 15573 2989 15673
rect 2589 15473 2989 15573
rect 2589 15373 2740 15473
rect 2840 15373 2989 15473
rect 2589 15273 2989 15373
rect 2589 15173 2740 15273
rect 2840 15173 2989 15273
rect 2589 15073 2989 15173
rect 2589 14973 2740 15073
rect 2840 14973 2989 15073
rect 2589 14707 2989 14973
rect 3089 17473 3489 17707
rect 3089 17373 3235 17473
rect 3335 17373 3489 17473
rect 3089 17273 3489 17373
rect 3089 17173 3235 17273
rect 3335 17173 3489 17273
rect 3089 17073 3489 17173
rect 3089 16973 3235 17073
rect 3335 16973 3489 17073
rect 3089 16873 3489 16973
rect 3089 16773 3235 16873
rect 3335 16773 3489 16873
rect 3089 16673 3489 16773
rect 3089 16573 3235 16673
rect 3335 16573 3489 16673
rect 3089 16473 3489 16573
rect 3089 16373 3235 16473
rect 3335 16373 3489 16473
rect 3089 16273 3489 16373
rect 3089 16173 3235 16273
rect 3335 16173 3489 16273
rect 3089 16073 3489 16173
rect 3089 15973 3235 16073
rect 3335 15973 3489 16073
rect 3089 15873 3489 15973
rect 3089 15773 3235 15873
rect 3335 15773 3489 15873
rect 3089 15673 3489 15773
rect 3089 15573 3235 15673
rect 3335 15573 3489 15673
rect 3089 15473 3489 15573
rect 3089 15373 3235 15473
rect 3335 15373 3489 15473
rect 3089 15273 3489 15373
rect 3089 15173 3235 15273
rect 3335 15173 3489 15273
rect 3089 15073 3489 15173
rect 3089 14973 3235 15073
rect 3335 14973 3489 15073
rect 3089 14707 3489 14973
rect 3589 17473 3989 17707
rect 3589 17373 3740 17473
rect 3840 17373 3989 17473
rect 3589 17273 3989 17373
rect 3589 17173 3740 17273
rect 3840 17173 3989 17273
rect 3589 17073 3989 17173
rect 3589 16973 3740 17073
rect 3840 16973 3989 17073
rect 3589 16873 3989 16973
rect 3589 16773 3740 16873
rect 3840 16773 3989 16873
rect 3589 16673 3989 16773
rect 3589 16573 3740 16673
rect 3840 16573 3989 16673
rect 3589 16473 3989 16573
rect 3589 16373 3740 16473
rect 3840 16373 3989 16473
rect 3589 16273 3989 16373
rect 3589 16173 3740 16273
rect 3840 16173 3989 16273
rect 3589 16073 3989 16173
rect 3589 15973 3740 16073
rect 3840 15973 3989 16073
rect 3589 15873 3989 15973
rect 3589 15773 3740 15873
rect 3840 15773 3989 15873
rect 3589 15673 3989 15773
rect 3589 15573 3740 15673
rect 3840 15573 3989 15673
rect 3589 15473 3989 15573
rect 3589 15373 3740 15473
rect 3840 15373 3989 15473
rect 3589 15273 3989 15373
rect 3589 15173 3740 15273
rect 3840 15173 3989 15273
rect 3589 15073 3989 15173
rect 3589 14973 3740 15073
rect 3840 14973 3989 15073
rect 3589 14707 3989 14973
rect 4089 17473 4489 17707
rect 4089 17373 4235 17473
rect 4335 17373 4489 17473
rect 4089 17273 4489 17373
rect 4089 17173 4235 17273
rect 4335 17173 4489 17273
rect 4089 17073 4489 17173
rect 4089 16973 4235 17073
rect 4335 16973 4489 17073
rect 4089 16873 4489 16973
rect 4089 16773 4235 16873
rect 4335 16773 4489 16873
rect 4089 16673 4489 16773
rect 4089 16573 4235 16673
rect 4335 16573 4489 16673
rect 4089 16473 4489 16573
rect 4089 16373 4235 16473
rect 4335 16373 4489 16473
rect 4089 16273 4489 16373
rect 4089 16173 4235 16273
rect 4335 16173 4489 16273
rect 4089 16073 4489 16173
rect 4089 15973 4235 16073
rect 4335 15973 4489 16073
rect 4089 15873 4489 15973
rect 4089 15773 4235 15873
rect 4335 15773 4489 15873
rect 4089 15673 4489 15773
rect 4089 15573 4235 15673
rect 4335 15573 4489 15673
rect 4089 15473 4489 15573
rect 4089 15373 4235 15473
rect 4335 15373 4489 15473
rect 4089 15273 4489 15373
rect 4089 15173 4235 15273
rect 4335 15173 4489 15273
rect 4089 15073 4489 15173
rect 4089 14973 4235 15073
rect 4335 14973 4489 15073
rect 4089 14707 4489 14973
rect 4589 17473 4989 17707
rect 4589 17373 4740 17473
rect 4840 17373 4989 17473
rect 4589 17273 4989 17373
rect 4589 17173 4740 17273
rect 4840 17173 4989 17273
rect 4589 17073 4989 17173
rect 4589 16973 4740 17073
rect 4840 16973 4989 17073
rect 4589 16873 4989 16973
rect 4589 16773 4740 16873
rect 4840 16773 4989 16873
rect 4589 16673 4989 16773
rect 4589 16573 4740 16673
rect 4840 16573 4989 16673
rect 4589 16473 4989 16573
rect 4589 16373 4740 16473
rect 4840 16373 4989 16473
rect 4589 16273 4989 16373
rect 4589 16173 4740 16273
rect 4840 16173 4989 16273
rect 4589 16073 4989 16173
rect 4589 15973 4740 16073
rect 4840 15973 4989 16073
rect 4589 15873 4989 15973
rect 4589 15773 4740 15873
rect 4840 15773 4989 15873
rect 4589 15673 4989 15773
rect 4589 15573 4740 15673
rect 4840 15573 4989 15673
rect 4589 15473 4989 15573
rect 4589 15373 4740 15473
rect 4840 15373 4989 15473
rect 4589 15273 4989 15373
rect 4589 15173 4740 15273
rect 4840 15173 4989 15273
rect 4589 15073 4989 15173
rect 4589 14973 4740 15073
rect 4840 14973 4989 15073
rect 4589 14707 4989 14973
rect 5089 17473 5489 17707
rect 5089 17373 5235 17473
rect 5335 17373 5489 17473
rect 5089 17273 5489 17373
rect 5089 17173 5235 17273
rect 5335 17173 5489 17273
rect 5089 17073 5489 17173
rect 5089 16973 5235 17073
rect 5335 16973 5489 17073
rect 5089 16873 5489 16973
rect 5089 16773 5235 16873
rect 5335 16773 5489 16873
rect 5089 16673 5489 16773
rect 5089 16573 5235 16673
rect 5335 16573 5489 16673
rect 5089 16473 5489 16573
rect 5089 16373 5235 16473
rect 5335 16373 5489 16473
rect 5089 16273 5489 16373
rect 5089 16173 5235 16273
rect 5335 16173 5489 16273
rect 5089 16073 5489 16173
rect 5089 15973 5235 16073
rect 5335 15973 5489 16073
rect 5089 15873 5489 15973
rect 5089 15773 5235 15873
rect 5335 15773 5489 15873
rect 5089 15673 5489 15773
rect 5089 15573 5235 15673
rect 5335 15573 5489 15673
rect 5089 15473 5489 15573
rect 5089 15373 5235 15473
rect 5335 15373 5489 15473
rect 5089 15273 5489 15373
rect 5089 15173 5235 15273
rect 5335 15173 5489 15273
rect 5089 15073 5489 15173
rect 5089 14973 5235 15073
rect 5335 14973 5489 15073
rect 5089 14707 5489 14973
rect 5589 17473 5989 17707
rect 5589 17373 5740 17473
rect 5840 17373 5989 17473
rect 5589 17273 5989 17373
rect 5589 17173 5740 17273
rect 5840 17173 5989 17273
rect 5589 17073 5989 17173
rect 5589 16973 5740 17073
rect 5840 16973 5989 17073
rect 5589 16873 5989 16973
rect 5589 16773 5740 16873
rect 5840 16773 5989 16873
rect 5589 16673 5989 16773
rect 5589 16573 5740 16673
rect 5840 16573 5989 16673
rect 5589 16473 5989 16573
rect 5589 16373 5740 16473
rect 5840 16373 5989 16473
rect 5589 16273 5989 16373
rect 5589 16173 5740 16273
rect 5840 16173 5989 16273
rect 5589 16073 5989 16173
rect 5589 15973 5740 16073
rect 5840 15973 5989 16073
rect 5589 15873 5989 15973
rect 5589 15773 5740 15873
rect 5840 15773 5989 15873
rect 5589 15673 5989 15773
rect 5589 15573 5740 15673
rect 5840 15573 5989 15673
rect 5589 15473 5989 15573
rect 5589 15373 5740 15473
rect 5840 15373 5989 15473
rect 5589 15273 5989 15373
rect 5589 15173 5740 15273
rect 5840 15173 5989 15273
rect 5589 15073 5989 15173
rect 5589 14973 5740 15073
rect 5840 14973 5989 15073
rect 5589 14707 5989 14973
rect 6089 17473 6489 17707
rect 6089 17373 6235 17473
rect 6335 17373 6489 17473
rect 6089 17273 6489 17373
rect 6089 17173 6235 17273
rect 6335 17173 6489 17273
rect 6089 17073 6489 17173
rect 6089 16973 6235 17073
rect 6335 16973 6489 17073
rect 6089 16873 6489 16973
rect 6089 16773 6235 16873
rect 6335 16773 6489 16873
rect 6089 16673 6489 16773
rect 6089 16573 6235 16673
rect 6335 16573 6489 16673
rect 6089 16473 6489 16573
rect 6089 16373 6235 16473
rect 6335 16373 6489 16473
rect 6089 16273 6489 16373
rect 6089 16173 6235 16273
rect 6335 16173 6489 16273
rect 6089 16073 6489 16173
rect 6089 15973 6235 16073
rect 6335 15973 6489 16073
rect 6089 15873 6489 15973
rect 6089 15773 6235 15873
rect 6335 15773 6489 15873
rect 6089 15673 6489 15773
rect 6089 15573 6235 15673
rect 6335 15573 6489 15673
rect 6089 15473 6489 15573
rect 6089 15373 6235 15473
rect 6335 15373 6489 15473
rect 6089 15273 6489 15373
rect 6089 15173 6235 15273
rect 6335 15173 6489 15273
rect 6089 15073 6489 15173
rect 6089 14973 6235 15073
rect 6335 14973 6489 15073
rect 6089 14707 6489 14973
rect 6589 17473 6989 17707
rect 6589 17373 6740 17473
rect 6840 17373 6989 17473
rect 6589 17273 6989 17373
rect 6589 17173 6740 17273
rect 6840 17173 6989 17273
rect 6589 17073 6989 17173
rect 6589 16973 6740 17073
rect 6840 16973 6989 17073
rect 6589 16873 6989 16973
rect 6589 16773 6740 16873
rect 6840 16773 6989 16873
rect 6589 16673 6989 16773
rect 6589 16573 6740 16673
rect 6840 16573 6989 16673
rect 6589 16473 6989 16573
rect 6589 16373 6740 16473
rect 6840 16373 6989 16473
rect 6589 16273 6989 16373
rect 6589 16173 6740 16273
rect 6840 16173 6989 16273
rect 6589 16073 6989 16173
rect 6589 15973 6740 16073
rect 6840 15973 6989 16073
rect 6589 15873 6989 15973
rect 6589 15773 6740 15873
rect 6840 15773 6989 15873
rect 6589 15673 6989 15773
rect 6589 15573 6740 15673
rect 6840 15573 6989 15673
rect 6589 15473 6989 15573
rect 6589 15373 6740 15473
rect 6840 15373 6989 15473
rect 6589 15273 6989 15373
rect 6589 15173 6740 15273
rect 6840 15173 6989 15273
rect 6589 15073 6989 15173
rect 6589 14973 6740 15073
rect 6840 14973 6989 15073
rect 6589 14707 6989 14973
rect 7089 17473 7489 17707
rect 7089 17373 7235 17473
rect 7335 17373 7489 17473
rect 7089 17273 7489 17373
rect 7089 17173 7235 17273
rect 7335 17173 7489 17273
rect 7089 17073 7489 17173
rect 7089 16973 7235 17073
rect 7335 16973 7489 17073
rect 7089 16873 7489 16973
rect 7089 16773 7235 16873
rect 7335 16773 7489 16873
rect 7089 16673 7489 16773
rect 7089 16573 7235 16673
rect 7335 16573 7489 16673
rect 7089 16473 7489 16573
rect 7089 16373 7235 16473
rect 7335 16373 7489 16473
rect 7089 16273 7489 16373
rect 7089 16173 7235 16273
rect 7335 16173 7489 16273
rect 7089 16073 7489 16173
rect 7089 15973 7235 16073
rect 7335 15973 7489 16073
rect 7089 15873 7489 15973
rect 7089 15773 7235 15873
rect 7335 15773 7489 15873
rect 7089 15673 7489 15773
rect 7089 15573 7235 15673
rect 7335 15573 7489 15673
rect 7089 15473 7489 15573
rect 7089 15373 7235 15473
rect 7335 15373 7489 15473
rect 7089 15273 7489 15373
rect 7089 15173 7235 15273
rect 7335 15173 7489 15273
rect 7089 15073 7489 15173
rect 7089 14973 7235 15073
rect 7335 14973 7489 15073
rect 7089 14707 7489 14973
rect 7589 17473 7989 17707
rect 7589 17373 7740 17473
rect 7840 17373 7989 17473
rect 7589 17273 7989 17373
rect 7589 17173 7740 17273
rect 7840 17173 7989 17273
rect 7589 17073 7989 17173
rect 7589 16973 7740 17073
rect 7840 16973 7989 17073
rect 7589 16873 7989 16973
rect 7589 16773 7740 16873
rect 7840 16773 7989 16873
rect 7589 16673 7989 16773
rect 7589 16573 7740 16673
rect 7840 16573 7989 16673
rect 7589 16473 7989 16573
rect 7589 16373 7740 16473
rect 7840 16373 7989 16473
rect 7589 16273 7989 16373
rect 7589 16173 7740 16273
rect 7840 16173 7989 16273
rect 7589 16073 7989 16173
rect 7589 15973 7740 16073
rect 7840 15973 7989 16073
rect 7589 15873 7989 15973
rect 7589 15773 7740 15873
rect 7840 15773 7989 15873
rect 7589 15673 7989 15773
rect 7589 15573 7740 15673
rect 7840 15573 7989 15673
rect 7589 15473 7989 15573
rect 7589 15373 7740 15473
rect 7840 15373 7989 15473
rect 7589 15273 7989 15373
rect 7589 15173 7740 15273
rect 7840 15173 7989 15273
rect 7589 15073 7989 15173
rect 7589 14973 7740 15073
rect 7840 14973 7989 15073
rect 7589 14707 7989 14973
rect 8089 17473 8489 17707
rect 8089 17373 8235 17473
rect 8335 17373 8489 17473
rect 8089 17273 8489 17373
rect 8089 17173 8235 17273
rect 8335 17173 8489 17273
rect 8089 17073 8489 17173
rect 8089 16973 8235 17073
rect 8335 16973 8489 17073
rect 8089 16873 8489 16973
rect 8089 16773 8235 16873
rect 8335 16773 8489 16873
rect 8089 16673 8489 16773
rect 8089 16573 8235 16673
rect 8335 16573 8489 16673
rect 8089 16473 8489 16573
rect 8089 16373 8235 16473
rect 8335 16373 8489 16473
rect 8089 16273 8489 16373
rect 8089 16173 8235 16273
rect 8335 16173 8489 16273
rect 8089 16073 8489 16173
rect 8089 15973 8235 16073
rect 8335 15973 8489 16073
rect 8089 15873 8489 15973
rect 8089 15773 8235 15873
rect 8335 15773 8489 15873
rect 8089 15673 8489 15773
rect 8089 15573 8235 15673
rect 8335 15573 8489 15673
rect 8089 15473 8489 15573
rect 8089 15373 8235 15473
rect 8335 15373 8489 15473
rect 8089 15273 8489 15373
rect 8089 15173 8235 15273
rect 8335 15173 8489 15273
rect 8089 15073 8489 15173
rect 8089 14973 8235 15073
rect 8335 14973 8489 15073
rect 8089 14707 8489 14973
rect 8589 17473 8989 17707
rect 8589 17373 8740 17473
rect 8840 17373 8989 17473
rect 8589 17273 8989 17373
rect 8589 17173 8740 17273
rect 8840 17173 8989 17273
rect 8589 17073 8989 17173
rect 8589 16973 8740 17073
rect 8840 16973 8989 17073
rect 8589 16873 8989 16973
rect 8589 16773 8740 16873
rect 8840 16773 8989 16873
rect 8589 16673 8989 16773
rect 8589 16573 8740 16673
rect 8840 16573 8989 16673
rect 8589 16473 8989 16573
rect 8589 16373 8740 16473
rect 8840 16373 8989 16473
rect 8589 16273 8989 16373
rect 8589 16173 8740 16273
rect 8840 16173 8989 16273
rect 8589 16073 8989 16173
rect 8589 15973 8740 16073
rect 8840 15973 8989 16073
rect 8589 15873 8989 15973
rect 8589 15773 8740 15873
rect 8840 15773 8989 15873
rect 8589 15673 8989 15773
rect 8589 15573 8740 15673
rect 8840 15573 8989 15673
rect 8589 15473 8989 15573
rect 8589 15373 8740 15473
rect 8840 15373 8989 15473
rect 8589 15273 8989 15373
rect 8589 15173 8740 15273
rect 8840 15173 8989 15273
rect 8589 15073 8989 15173
rect 8589 14973 8740 15073
rect 8840 14973 8989 15073
rect 8589 14707 8989 14973
rect 9089 17473 9489 17707
rect 9089 17373 9235 17473
rect 9335 17373 9489 17473
rect 9089 17273 9489 17373
rect 9089 17173 9235 17273
rect 9335 17173 9489 17273
rect 9089 17073 9489 17173
rect 9089 16973 9235 17073
rect 9335 16973 9489 17073
rect 9089 16873 9489 16973
rect 9089 16773 9235 16873
rect 9335 16773 9489 16873
rect 9089 16673 9489 16773
rect 9089 16573 9235 16673
rect 9335 16573 9489 16673
rect 9089 16473 9489 16573
rect 9089 16373 9235 16473
rect 9335 16373 9489 16473
rect 9089 16273 9489 16373
rect 9089 16173 9235 16273
rect 9335 16173 9489 16273
rect 9089 16073 9489 16173
rect 9089 15973 9235 16073
rect 9335 15973 9489 16073
rect 9089 15873 9489 15973
rect 9089 15773 9235 15873
rect 9335 15773 9489 15873
rect 9089 15673 9489 15773
rect 9089 15573 9235 15673
rect 9335 15573 9489 15673
rect 9089 15473 9489 15573
rect 9089 15373 9235 15473
rect 9335 15373 9489 15473
rect 9089 15273 9489 15373
rect 9089 15173 9235 15273
rect 9335 15173 9489 15273
rect 9089 15073 9489 15173
rect 9089 14973 9235 15073
rect 9335 14973 9489 15073
rect 9089 14707 9489 14973
rect 9589 17473 10031 17707
rect 9589 17373 9740 17473
rect 9840 17373 10031 17473
rect 9589 17273 10031 17373
rect 9589 17173 9740 17273
rect 9840 17173 10031 17273
rect 9589 17073 10031 17173
rect 9589 16973 9740 17073
rect 9840 16973 10031 17073
rect 9589 16873 10031 16973
rect 9589 16773 9740 16873
rect 9840 16773 10031 16873
rect 9589 16673 10031 16773
rect 9589 16573 9740 16673
rect 9840 16573 10031 16673
rect 9589 16473 10031 16573
rect 9589 16373 9740 16473
rect 9840 16373 10031 16473
rect 9589 16273 10031 16373
rect 9589 16173 9740 16273
rect 9840 16173 10031 16273
rect 9589 16073 10031 16173
rect 9589 15973 9740 16073
rect 9840 15973 10031 16073
rect 9589 15873 10031 15973
rect 9589 15773 9740 15873
rect 9840 15773 10031 15873
rect 9589 15673 10031 15773
rect 9589 15573 9740 15673
rect 9840 15573 10031 15673
rect 9589 15473 10031 15573
rect 9589 15373 9740 15473
rect 9840 15373 10031 15473
rect 9589 15273 10031 15373
rect 9589 15173 9740 15273
rect 9840 15173 10031 15273
rect 9589 15073 10031 15173
rect 9589 14973 9740 15073
rect 9840 14973 10031 15073
rect 9589 14707 10031 14973
rect -433 11746 9 12012
rect -433 11646 -242 11746
rect -142 11646 9 11746
rect -433 11546 9 11646
rect -433 11446 -242 11546
rect -142 11446 9 11546
rect -433 11346 9 11446
rect -433 11246 -242 11346
rect -142 11246 9 11346
rect -433 11146 9 11246
rect -433 11046 -242 11146
rect -142 11046 9 11146
rect -433 10946 9 11046
rect -433 10846 -242 10946
rect -142 10846 9 10946
rect -433 10746 9 10846
rect -433 10646 -242 10746
rect -142 10646 9 10746
rect -433 10546 9 10646
rect -433 10446 -242 10546
rect -142 10446 9 10546
rect -433 10346 9 10446
rect -433 10246 -242 10346
rect -142 10246 9 10346
rect -433 10146 9 10246
rect -433 10046 -242 10146
rect -142 10046 9 10146
rect -433 9946 9 10046
rect -433 9846 -242 9946
rect -142 9846 9 9946
rect -433 9746 9 9846
rect -433 9646 -242 9746
rect -142 9646 9 9746
rect -433 9546 9 9646
rect -433 9446 -242 9546
rect -142 9446 9 9546
rect -433 9346 9 9446
rect -433 9246 -242 9346
rect -142 9246 9 9346
rect -433 9012 9 9246
rect 109 11746 509 12012
rect 109 11646 263 11746
rect 363 11646 509 11746
rect 109 11546 509 11646
rect 109 11446 263 11546
rect 363 11446 509 11546
rect 109 11346 509 11446
rect 109 11246 263 11346
rect 363 11246 509 11346
rect 109 11146 509 11246
rect 109 11046 263 11146
rect 363 11046 509 11146
rect 109 10946 509 11046
rect 109 10846 263 10946
rect 363 10846 509 10946
rect 109 10746 509 10846
rect 109 10646 263 10746
rect 363 10646 509 10746
rect 109 10546 509 10646
rect 109 10446 263 10546
rect 363 10446 509 10546
rect 109 10346 509 10446
rect 109 10246 263 10346
rect 363 10246 509 10346
rect 109 10146 509 10246
rect 109 10046 263 10146
rect 363 10046 509 10146
rect 109 9946 509 10046
rect 109 9846 263 9946
rect 363 9846 509 9946
rect 109 9746 509 9846
rect 109 9646 263 9746
rect 363 9646 509 9746
rect 109 9546 509 9646
rect 109 9446 263 9546
rect 363 9446 509 9546
rect 109 9346 509 9446
rect 109 9246 263 9346
rect 363 9246 509 9346
rect 109 9012 509 9246
rect 609 11746 1009 12012
rect 609 11646 758 11746
rect 858 11646 1009 11746
rect 609 11546 1009 11646
rect 609 11446 758 11546
rect 858 11446 1009 11546
rect 609 11346 1009 11446
rect 609 11246 758 11346
rect 858 11246 1009 11346
rect 609 11146 1009 11246
rect 609 11046 758 11146
rect 858 11046 1009 11146
rect 609 10946 1009 11046
rect 609 10846 758 10946
rect 858 10846 1009 10946
rect 609 10746 1009 10846
rect 609 10646 758 10746
rect 858 10646 1009 10746
rect 609 10546 1009 10646
rect 609 10446 758 10546
rect 858 10446 1009 10546
rect 609 10346 1009 10446
rect 609 10246 758 10346
rect 858 10246 1009 10346
rect 609 10146 1009 10246
rect 609 10046 758 10146
rect 858 10046 1009 10146
rect 609 9946 1009 10046
rect 609 9846 758 9946
rect 858 9846 1009 9946
rect 609 9746 1009 9846
rect 609 9646 758 9746
rect 858 9646 1009 9746
rect 609 9546 1009 9646
rect 609 9446 758 9546
rect 858 9446 1009 9546
rect 609 9346 1009 9446
rect 609 9246 758 9346
rect 858 9246 1009 9346
rect 609 9012 1009 9246
rect 1109 11746 1509 12012
rect 1109 11646 1263 11746
rect 1363 11646 1509 11746
rect 1109 11546 1509 11646
rect 1109 11446 1263 11546
rect 1363 11446 1509 11546
rect 1109 11346 1509 11446
rect 1109 11246 1263 11346
rect 1363 11246 1509 11346
rect 1109 11146 1509 11246
rect 1109 11046 1263 11146
rect 1363 11046 1509 11146
rect 1109 10946 1509 11046
rect 1109 10846 1263 10946
rect 1363 10846 1509 10946
rect 1109 10746 1509 10846
rect 1109 10646 1263 10746
rect 1363 10646 1509 10746
rect 1109 10546 1509 10646
rect 1109 10446 1263 10546
rect 1363 10446 1509 10546
rect 1109 10346 1509 10446
rect 1109 10246 1263 10346
rect 1363 10246 1509 10346
rect 1109 10146 1509 10246
rect 1109 10046 1263 10146
rect 1363 10046 1509 10146
rect 1109 9946 1509 10046
rect 1109 9846 1263 9946
rect 1363 9846 1509 9946
rect 1109 9746 1509 9846
rect 1109 9646 1263 9746
rect 1363 9646 1509 9746
rect 1109 9546 1509 9646
rect 1109 9446 1263 9546
rect 1363 9446 1509 9546
rect 1109 9346 1509 9446
rect 1109 9246 1263 9346
rect 1363 9246 1509 9346
rect 1109 9012 1509 9246
rect 1609 11746 2009 12012
rect 1609 11646 1758 11746
rect 1858 11646 2009 11746
rect 1609 11546 2009 11646
rect 1609 11446 1758 11546
rect 1858 11446 2009 11546
rect 1609 11346 2009 11446
rect 1609 11246 1758 11346
rect 1858 11246 2009 11346
rect 1609 11146 2009 11246
rect 1609 11046 1758 11146
rect 1858 11046 2009 11146
rect 1609 10946 2009 11046
rect 1609 10846 1758 10946
rect 1858 10846 2009 10946
rect 1609 10746 2009 10846
rect 1609 10646 1758 10746
rect 1858 10646 2009 10746
rect 1609 10546 2009 10646
rect 1609 10446 1758 10546
rect 1858 10446 2009 10546
rect 1609 10346 2009 10446
rect 1609 10246 1758 10346
rect 1858 10246 2009 10346
rect 1609 10146 2009 10246
rect 1609 10046 1758 10146
rect 1858 10046 2009 10146
rect 1609 9946 2009 10046
rect 1609 9846 1758 9946
rect 1858 9846 2009 9946
rect 1609 9746 2009 9846
rect 1609 9646 1758 9746
rect 1858 9646 2009 9746
rect 1609 9546 2009 9646
rect 1609 9446 1758 9546
rect 1858 9446 2009 9546
rect 1609 9346 2009 9446
rect 1609 9246 1758 9346
rect 1858 9246 2009 9346
rect 1609 9012 2009 9246
rect 2109 11746 2509 12012
rect 2109 11646 2263 11746
rect 2363 11646 2509 11746
rect 2109 11546 2509 11646
rect 2109 11446 2263 11546
rect 2363 11446 2509 11546
rect 2109 11346 2509 11446
rect 2109 11246 2263 11346
rect 2363 11246 2509 11346
rect 2109 11146 2509 11246
rect 2109 11046 2263 11146
rect 2363 11046 2509 11146
rect 2109 10946 2509 11046
rect 2109 10846 2263 10946
rect 2363 10846 2509 10946
rect 2109 10746 2509 10846
rect 2109 10646 2263 10746
rect 2363 10646 2509 10746
rect 2109 10546 2509 10646
rect 2109 10446 2263 10546
rect 2363 10446 2509 10546
rect 2109 10346 2509 10446
rect 2109 10246 2263 10346
rect 2363 10246 2509 10346
rect 2109 10146 2509 10246
rect 2109 10046 2263 10146
rect 2363 10046 2509 10146
rect 2109 9946 2509 10046
rect 2109 9846 2263 9946
rect 2363 9846 2509 9946
rect 2109 9746 2509 9846
rect 2109 9646 2263 9746
rect 2363 9646 2509 9746
rect 2109 9546 2509 9646
rect 2109 9446 2263 9546
rect 2363 9446 2509 9546
rect 2109 9346 2509 9446
rect 2109 9246 2263 9346
rect 2363 9246 2509 9346
rect 2109 9012 2509 9246
rect 2609 11746 3009 12012
rect 2609 11646 2758 11746
rect 2858 11646 3009 11746
rect 2609 11546 3009 11646
rect 2609 11446 2758 11546
rect 2858 11446 3009 11546
rect 2609 11346 3009 11446
rect 2609 11246 2758 11346
rect 2858 11246 3009 11346
rect 2609 11146 3009 11246
rect 2609 11046 2758 11146
rect 2858 11046 3009 11146
rect 2609 10946 3009 11046
rect 2609 10846 2758 10946
rect 2858 10846 3009 10946
rect 2609 10746 3009 10846
rect 2609 10646 2758 10746
rect 2858 10646 3009 10746
rect 2609 10546 3009 10646
rect 2609 10446 2758 10546
rect 2858 10446 3009 10546
rect 2609 10346 3009 10446
rect 2609 10246 2758 10346
rect 2858 10246 3009 10346
rect 2609 10146 3009 10246
rect 2609 10046 2758 10146
rect 2858 10046 3009 10146
rect 2609 9946 3009 10046
rect 2609 9846 2758 9946
rect 2858 9846 3009 9946
rect 2609 9746 3009 9846
rect 2609 9646 2758 9746
rect 2858 9646 3009 9746
rect 2609 9546 3009 9646
rect 2609 9446 2758 9546
rect 2858 9446 3009 9546
rect 2609 9346 3009 9446
rect 2609 9246 2758 9346
rect 2858 9246 3009 9346
rect 2609 9012 3009 9246
rect 3109 11746 3509 12012
rect 3109 11646 3263 11746
rect 3363 11646 3509 11746
rect 3109 11546 3509 11646
rect 3109 11446 3263 11546
rect 3363 11446 3509 11546
rect 3109 11346 3509 11446
rect 3109 11246 3263 11346
rect 3363 11246 3509 11346
rect 3109 11146 3509 11246
rect 3109 11046 3263 11146
rect 3363 11046 3509 11146
rect 3109 10946 3509 11046
rect 3109 10846 3263 10946
rect 3363 10846 3509 10946
rect 3109 10746 3509 10846
rect 3109 10646 3263 10746
rect 3363 10646 3509 10746
rect 3109 10546 3509 10646
rect 3109 10446 3263 10546
rect 3363 10446 3509 10546
rect 3109 10346 3509 10446
rect 3109 10246 3263 10346
rect 3363 10246 3509 10346
rect 3109 10146 3509 10246
rect 3109 10046 3263 10146
rect 3363 10046 3509 10146
rect 3109 9946 3509 10046
rect 3109 9846 3263 9946
rect 3363 9846 3509 9946
rect 3109 9746 3509 9846
rect 3109 9646 3263 9746
rect 3363 9646 3509 9746
rect 3109 9546 3509 9646
rect 3109 9446 3263 9546
rect 3363 9446 3509 9546
rect 3109 9346 3509 9446
rect 3109 9246 3263 9346
rect 3363 9246 3509 9346
rect 3109 9012 3509 9246
rect 3609 11746 4009 12012
rect 3609 11646 3758 11746
rect 3858 11646 4009 11746
rect 3609 11546 4009 11646
rect 3609 11446 3758 11546
rect 3858 11446 4009 11546
rect 3609 11346 4009 11446
rect 3609 11246 3758 11346
rect 3858 11246 4009 11346
rect 3609 11146 4009 11246
rect 3609 11046 3758 11146
rect 3858 11046 4009 11146
rect 3609 10946 4009 11046
rect 3609 10846 3758 10946
rect 3858 10846 4009 10946
rect 3609 10746 4009 10846
rect 3609 10646 3758 10746
rect 3858 10646 4009 10746
rect 3609 10546 4009 10646
rect 3609 10446 3758 10546
rect 3858 10446 4009 10546
rect 3609 10346 4009 10446
rect 3609 10246 3758 10346
rect 3858 10246 4009 10346
rect 3609 10146 4009 10246
rect 3609 10046 3758 10146
rect 3858 10046 4009 10146
rect 3609 9946 4009 10046
rect 3609 9846 3758 9946
rect 3858 9846 4009 9946
rect 3609 9746 4009 9846
rect 3609 9646 3758 9746
rect 3858 9646 4009 9746
rect 3609 9546 4009 9646
rect 3609 9446 3758 9546
rect 3858 9446 4009 9546
rect 3609 9346 4009 9446
rect 3609 9246 3758 9346
rect 3858 9246 4009 9346
rect 3609 9012 4009 9246
rect 4109 11746 4509 12012
rect 4109 11646 4263 11746
rect 4363 11646 4509 11746
rect 4109 11546 4509 11646
rect 4109 11446 4263 11546
rect 4363 11446 4509 11546
rect 4109 11346 4509 11446
rect 4109 11246 4263 11346
rect 4363 11246 4509 11346
rect 4109 11146 4509 11246
rect 4109 11046 4263 11146
rect 4363 11046 4509 11146
rect 4109 10946 4509 11046
rect 4109 10846 4263 10946
rect 4363 10846 4509 10946
rect 4109 10746 4509 10846
rect 4109 10646 4263 10746
rect 4363 10646 4509 10746
rect 4109 10546 4509 10646
rect 4109 10446 4263 10546
rect 4363 10446 4509 10546
rect 4109 10346 4509 10446
rect 4109 10246 4263 10346
rect 4363 10246 4509 10346
rect 4109 10146 4509 10246
rect 4109 10046 4263 10146
rect 4363 10046 4509 10146
rect 4109 9946 4509 10046
rect 4109 9846 4263 9946
rect 4363 9846 4509 9946
rect 4109 9746 4509 9846
rect 4109 9646 4263 9746
rect 4363 9646 4509 9746
rect 4109 9546 4509 9646
rect 4109 9446 4263 9546
rect 4363 9446 4509 9546
rect 4109 9346 4509 9446
rect 4109 9246 4263 9346
rect 4363 9246 4509 9346
rect 4109 9012 4509 9246
rect 4609 11746 5009 12012
rect 4609 11646 4758 11746
rect 4858 11646 5009 11746
rect 4609 11546 5009 11646
rect 4609 11446 4758 11546
rect 4858 11446 5009 11546
rect 4609 11346 5009 11446
rect 4609 11246 4758 11346
rect 4858 11246 5009 11346
rect 4609 11146 5009 11246
rect 4609 11046 4758 11146
rect 4858 11046 5009 11146
rect 4609 10946 5009 11046
rect 4609 10846 4758 10946
rect 4858 10846 5009 10946
rect 4609 10746 5009 10846
rect 4609 10646 4758 10746
rect 4858 10646 5009 10746
rect 4609 10546 5009 10646
rect 4609 10446 4758 10546
rect 4858 10446 5009 10546
rect 4609 10346 5009 10446
rect 4609 10246 4758 10346
rect 4858 10246 5009 10346
rect 4609 10146 5009 10246
rect 4609 10046 4758 10146
rect 4858 10046 5009 10146
rect 4609 9946 5009 10046
rect 4609 9846 4758 9946
rect 4858 9846 5009 9946
rect 4609 9746 5009 9846
rect 4609 9646 4758 9746
rect 4858 9646 5009 9746
rect 4609 9546 5009 9646
rect 4609 9446 4758 9546
rect 4858 9446 5009 9546
rect 4609 9346 5009 9446
rect 4609 9246 4758 9346
rect 4858 9246 5009 9346
rect 4609 9012 5009 9246
rect 5109 11746 5509 12012
rect 5109 11646 5263 11746
rect 5363 11646 5509 11746
rect 5109 11546 5509 11646
rect 5109 11446 5263 11546
rect 5363 11446 5509 11546
rect 5109 11346 5509 11446
rect 5109 11246 5263 11346
rect 5363 11246 5509 11346
rect 5109 11146 5509 11246
rect 5109 11046 5263 11146
rect 5363 11046 5509 11146
rect 5109 10946 5509 11046
rect 5109 10846 5263 10946
rect 5363 10846 5509 10946
rect 5109 10746 5509 10846
rect 5109 10646 5263 10746
rect 5363 10646 5509 10746
rect 5109 10546 5509 10646
rect 5109 10446 5263 10546
rect 5363 10446 5509 10546
rect 5109 10346 5509 10446
rect 5109 10246 5263 10346
rect 5363 10246 5509 10346
rect 5109 10146 5509 10246
rect 5109 10046 5263 10146
rect 5363 10046 5509 10146
rect 5109 9946 5509 10046
rect 5109 9846 5263 9946
rect 5363 9846 5509 9946
rect 5109 9746 5509 9846
rect 5109 9646 5263 9746
rect 5363 9646 5509 9746
rect 5109 9546 5509 9646
rect 5109 9446 5263 9546
rect 5363 9446 5509 9546
rect 5109 9346 5509 9446
rect 5109 9246 5263 9346
rect 5363 9246 5509 9346
rect 5109 9012 5509 9246
rect 5609 11746 6009 12012
rect 5609 11646 5758 11746
rect 5858 11646 6009 11746
rect 5609 11546 6009 11646
rect 5609 11446 5758 11546
rect 5858 11446 6009 11546
rect 5609 11346 6009 11446
rect 5609 11246 5758 11346
rect 5858 11246 6009 11346
rect 5609 11146 6009 11246
rect 5609 11046 5758 11146
rect 5858 11046 6009 11146
rect 5609 10946 6009 11046
rect 5609 10846 5758 10946
rect 5858 10846 6009 10946
rect 5609 10746 6009 10846
rect 5609 10646 5758 10746
rect 5858 10646 6009 10746
rect 5609 10546 6009 10646
rect 5609 10446 5758 10546
rect 5858 10446 6009 10546
rect 5609 10346 6009 10446
rect 5609 10246 5758 10346
rect 5858 10246 6009 10346
rect 5609 10146 6009 10246
rect 5609 10046 5758 10146
rect 5858 10046 6009 10146
rect 5609 9946 6009 10046
rect 5609 9846 5758 9946
rect 5858 9846 6009 9946
rect 5609 9746 6009 9846
rect 5609 9646 5758 9746
rect 5858 9646 6009 9746
rect 5609 9546 6009 9646
rect 5609 9446 5758 9546
rect 5858 9446 6009 9546
rect 5609 9346 6009 9446
rect 5609 9246 5758 9346
rect 5858 9246 6009 9346
rect 5609 9012 6009 9246
rect 6109 11746 6509 12012
rect 6109 11646 6263 11746
rect 6363 11646 6509 11746
rect 6109 11546 6509 11646
rect 6109 11446 6263 11546
rect 6363 11446 6509 11546
rect 6109 11346 6509 11446
rect 6109 11246 6263 11346
rect 6363 11246 6509 11346
rect 6109 11146 6509 11246
rect 6109 11046 6263 11146
rect 6363 11046 6509 11146
rect 6109 10946 6509 11046
rect 6109 10846 6263 10946
rect 6363 10846 6509 10946
rect 6109 10746 6509 10846
rect 6109 10646 6263 10746
rect 6363 10646 6509 10746
rect 6109 10546 6509 10646
rect 6109 10446 6263 10546
rect 6363 10446 6509 10546
rect 6109 10346 6509 10446
rect 6109 10246 6263 10346
rect 6363 10246 6509 10346
rect 6109 10146 6509 10246
rect 6109 10046 6263 10146
rect 6363 10046 6509 10146
rect 6109 9946 6509 10046
rect 6109 9846 6263 9946
rect 6363 9846 6509 9946
rect 6109 9746 6509 9846
rect 6109 9646 6263 9746
rect 6363 9646 6509 9746
rect 6109 9546 6509 9646
rect 6109 9446 6263 9546
rect 6363 9446 6509 9546
rect 6109 9346 6509 9446
rect 6109 9246 6263 9346
rect 6363 9246 6509 9346
rect 6109 9012 6509 9246
rect 6609 11746 7009 12012
rect 6609 11646 6758 11746
rect 6858 11646 7009 11746
rect 6609 11546 7009 11646
rect 6609 11446 6758 11546
rect 6858 11446 7009 11546
rect 6609 11346 7009 11446
rect 6609 11246 6758 11346
rect 6858 11246 7009 11346
rect 6609 11146 7009 11246
rect 6609 11046 6758 11146
rect 6858 11046 7009 11146
rect 6609 10946 7009 11046
rect 6609 10846 6758 10946
rect 6858 10846 7009 10946
rect 6609 10746 7009 10846
rect 6609 10646 6758 10746
rect 6858 10646 7009 10746
rect 6609 10546 7009 10646
rect 6609 10446 6758 10546
rect 6858 10446 7009 10546
rect 6609 10346 7009 10446
rect 6609 10246 6758 10346
rect 6858 10246 7009 10346
rect 6609 10146 7009 10246
rect 6609 10046 6758 10146
rect 6858 10046 7009 10146
rect 6609 9946 7009 10046
rect 6609 9846 6758 9946
rect 6858 9846 7009 9946
rect 6609 9746 7009 9846
rect 6609 9646 6758 9746
rect 6858 9646 7009 9746
rect 6609 9546 7009 9646
rect 6609 9446 6758 9546
rect 6858 9446 7009 9546
rect 6609 9346 7009 9446
rect 6609 9246 6758 9346
rect 6858 9246 7009 9346
rect 6609 9012 7009 9246
rect 7109 11746 7509 12012
rect 7109 11646 7263 11746
rect 7363 11646 7509 11746
rect 7109 11546 7509 11646
rect 7109 11446 7263 11546
rect 7363 11446 7509 11546
rect 7109 11346 7509 11446
rect 7109 11246 7263 11346
rect 7363 11246 7509 11346
rect 7109 11146 7509 11246
rect 7109 11046 7263 11146
rect 7363 11046 7509 11146
rect 7109 10946 7509 11046
rect 7109 10846 7263 10946
rect 7363 10846 7509 10946
rect 7109 10746 7509 10846
rect 7109 10646 7263 10746
rect 7363 10646 7509 10746
rect 7109 10546 7509 10646
rect 7109 10446 7263 10546
rect 7363 10446 7509 10546
rect 7109 10346 7509 10446
rect 7109 10246 7263 10346
rect 7363 10246 7509 10346
rect 7109 10146 7509 10246
rect 7109 10046 7263 10146
rect 7363 10046 7509 10146
rect 7109 9946 7509 10046
rect 7109 9846 7263 9946
rect 7363 9846 7509 9946
rect 7109 9746 7509 9846
rect 7109 9646 7263 9746
rect 7363 9646 7509 9746
rect 7109 9546 7509 9646
rect 7109 9446 7263 9546
rect 7363 9446 7509 9546
rect 7109 9346 7509 9446
rect 7109 9246 7263 9346
rect 7363 9246 7509 9346
rect 7109 9012 7509 9246
rect 7609 11746 8009 12012
rect 7609 11646 7758 11746
rect 7858 11646 8009 11746
rect 7609 11546 8009 11646
rect 7609 11446 7758 11546
rect 7858 11446 8009 11546
rect 7609 11346 8009 11446
rect 7609 11246 7758 11346
rect 7858 11246 8009 11346
rect 7609 11146 8009 11246
rect 7609 11046 7758 11146
rect 7858 11046 8009 11146
rect 7609 10946 8009 11046
rect 7609 10846 7758 10946
rect 7858 10846 8009 10946
rect 7609 10746 8009 10846
rect 7609 10646 7758 10746
rect 7858 10646 8009 10746
rect 7609 10546 8009 10646
rect 7609 10446 7758 10546
rect 7858 10446 8009 10546
rect 7609 10346 8009 10446
rect 7609 10246 7758 10346
rect 7858 10246 8009 10346
rect 7609 10146 8009 10246
rect 7609 10046 7758 10146
rect 7858 10046 8009 10146
rect 7609 9946 8009 10046
rect 7609 9846 7758 9946
rect 7858 9846 8009 9946
rect 7609 9746 8009 9846
rect 7609 9646 7758 9746
rect 7858 9646 8009 9746
rect 7609 9546 8009 9646
rect 7609 9446 7758 9546
rect 7858 9446 8009 9546
rect 7609 9346 8009 9446
rect 7609 9246 7758 9346
rect 7858 9246 8009 9346
rect 7609 9012 8009 9246
rect 8109 11746 8509 12012
rect 8109 11646 8263 11746
rect 8363 11646 8509 11746
rect 8109 11546 8509 11646
rect 8109 11446 8263 11546
rect 8363 11446 8509 11546
rect 8109 11346 8509 11446
rect 8109 11246 8263 11346
rect 8363 11246 8509 11346
rect 8109 11146 8509 11246
rect 8109 11046 8263 11146
rect 8363 11046 8509 11146
rect 8109 10946 8509 11046
rect 8109 10846 8263 10946
rect 8363 10846 8509 10946
rect 8109 10746 8509 10846
rect 8109 10646 8263 10746
rect 8363 10646 8509 10746
rect 8109 10546 8509 10646
rect 8109 10446 8263 10546
rect 8363 10446 8509 10546
rect 8109 10346 8509 10446
rect 8109 10246 8263 10346
rect 8363 10246 8509 10346
rect 8109 10146 8509 10246
rect 8109 10046 8263 10146
rect 8363 10046 8509 10146
rect 8109 9946 8509 10046
rect 8109 9846 8263 9946
rect 8363 9846 8509 9946
rect 8109 9746 8509 9846
rect 8109 9646 8263 9746
rect 8363 9646 8509 9746
rect 8109 9546 8509 9646
rect 8109 9446 8263 9546
rect 8363 9446 8509 9546
rect 8109 9346 8509 9446
rect 8109 9246 8263 9346
rect 8363 9246 8509 9346
rect 8109 9012 8509 9246
rect 8609 11746 9009 12012
rect 8609 11646 8758 11746
rect 8858 11646 9009 11746
rect 8609 11546 9009 11646
rect 8609 11446 8758 11546
rect 8858 11446 9009 11546
rect 8609 11346 9009 11446
rect 8609 11246 8758 11346
rect 8858 11246 9009 11346
rect 8609 11146 9009 11246
rect 8609 11046 8758 11146
rect 8858 11046 9009 11146
rect 8609 10946 9009 11046
rect 8609 10846 8758 10946
rect 8858 10846 9009 10946
rect 8609 10746 9009 10846
rect 8609 10646 8758 10746
rect 8858 10646 9009 10746
rect 8609 10546 9009 10646
rect 8609 10446 8758 10546
rect 8858 10446 9009 10546
rect 8609 10346 9009 10446
rect 8609 10246 8758 10346
rect 8858 10246 9009 10346
rect 8609 10146 9009 10246
rect 8609 10046 8758 10146
rect 8858 10046 9009 10146
rect 8609 9946 9009 10046
rect 8609 9846 8758 9946
rect 8858 9846 9009 9946
rect 8609 9746 9009 9846
rect 8609 9646 8758 9746
rect 8858 9646 9009 9746
rect 8609 9546 9009 9646
rect 8609 9446 8758 9546
rect 8858 9446 9009 9546
rect 8609 9346 9009 9446
rect 8609 9246 8758 9346
rect 8858 9246 9009 9346
rect 8609 9012 9009 9246
rect 9109 11746 9509 12012
rect 9109 11646 9263 11746
rect 9363 11646 9509 11746
rect 9109 11546 9509 11646
rect 9109 11446 9263 11546
rect 9363 11446 9509 11546
rect 9109 11346 9509 11446
rect 9109 11246 9263 11346
rect 9363 11246 9509 11346
rect 9109 11146 9509 11246
rect 9109 11046 9263 11146
rect 9363 11046 9509 11146
rect 9109 10946 9509 11046
rect 9109 10846 9263 10946
rect 9363 10846 9509 10946
rect 9109 10746 9509 10846
rect 9109 10646 9263 10746
rect 9363 10646 9509 10746
rect 9109 10546 9509 10646
rect 9109 10446 9263 10546
rect 9363 10446 9509 10546
rect 9109 10346 9509 10446
rect 9109 10246 9263 10346
rect 9363 10246 9509 10346
rect 9109 10146 9509 10246
rect 9109 10046 9263 10146
rect 9363 10046 9509 10146
rect 9109 9946 9509 10046
rect 9109 9846 9263 9946
rect 9363 9846 9509 9946
rect 9109 9746 9509 9846
rect 9109 9646 9263 9746
rect 9363 9646 9509 9746
rect 9109 9546 9509 9646
rect 9109 9446 9263 9546
rect 9363 9446 9509 9546
rect 9109 9346 9509 9446
rect 9109 9246 9263 9346
rect 9363 9246 9509 9346
rect 9109 9012 9509 9246
rect 9609 11742 10067 12012
rect 9609 11642 9782 11742
rect 9882 11642 10067 11742
rect 9609 11542 10067 11642
rect 9609 11442 9782 11542
rect 9882 11442 10067 11542
rect 9609 11342 10067 11442
rect 9609 11242 9782 11342
rect 9882 11242 10067 11342
rect 9609 11142 10067 11242
rect 9609 11042 9782 11142
rect 9882 11042 10067 11142
rect 9609 10942 10067 11042
rect 9609 10842 9782 10942
rect 9882 10842 10067 10942
rect 9609 10742 10067 10842
rect 9609 10642 9782 10742
rect 9882 10642 10067 10742
rect 9609 10542 10067 10642
rect 9609 10442 9782 10542
rect 9882 10442 10067 10542
rect 9609 10342 10067 10442
rect 9609 10242 9782 10342
rect 9882 10242 10067 10342
rect 9609 10142 10067 10242
rect 9609 10042 9782 10142
rect 9882 10042 10067 10142
rect 9609 9942 10067 10042
rect 9609 9842 9782 9942
rect 9882 9842 10067 9942
rect 9609 9742 10067 9842
rect 9609 9642 9782 9742
rect 9882 9642 10067 9742
rect 9609 9542 10067 9642
rect 9609 9442 9782 9542
rect 9882 9442 10067 9542
rect 9609 9342 10067 9442
rect 9609 9242 9782 9342
rect 9882 9242 10067 9342
rect 9609 9012 10067 9242
<< ndiffc >>
rect -104 6757 16 6857
rect -104 6557 16 6657
rect -104 6357 16 6457
rect -104 6157 16 6257
rect -104 5957 16 6057
rect 242 6757 362 6857
rect 242 6557 362 6657
rect 242 6357 362 6457
rect 242 6157 362 6257
rect 242 5957 362 6057
rect 648 6757 768 6857
rect 648 6557 768 6657
rect 648 6357 768 6457
rect 648 6157 768 6257
rect 648 5957 768 6057
rect 1018 6757 1138 6857
rect 1018 6557 1138 6657
rect 1018 6357 1138 6457
rect 1018 6157 1138 6257
rect 1018 5957 1138 6057
rect 1424 6757 1544 6857
rect 1424 6557 1544 6657
rect 1424 6357 1544 6457
rect 1424 6157 1544 6257
rect 1424 5957 1544 6057
rect 1770 6757 1890 6857
rect 1770 6557 1890 6657
rect 1770 6357 1890 6457
rect 1770 6157 1890 6257
rect 1770 5957 1890 6057
<< pdiffc >>
rect -284 17377 -184 17477
rect -284 17177 -184 17277
rect -284 16977 -184 17077
rect -284 16777 -184 16877
rect -284 16577 -184 16677
rect -284 16377 -184 16477
rect -284 16177 -184 16277
rect -284 15977 -184 16077
rect -284 15777 -184 15877
rect -284 15577 -184 15677
rect -284 15377 -184 15477
rect -284 15177 -184 15277
rect -284 14977 -184 15077
rect 235 17373 335 17473
rect 235 17173 335 17273
rect 235 16973 335 17073
rect 235 16773 335 16873
rect 235 16573 335 16673
rect 235 16373 335 16473
rect 235 16173 335 16273
rect 235 15973 335 16073
rect 235 15773 335 15873
rect 235 15573 335 15673
rect 235 15373 335 15473
rect 235 15173 335 15273
rect 235 14973 335 15073
rect 740 17373 840 17473
rect 740 17173 840 17273
rect 740 16973 840 17073
rect 740 16773 840 16873
rect 740 16573 840 16673
rect 740 16373 840 16473
rect 740 16173 840 16273
rect 740 15973 840 16073
rect 740 15773 840 15873
rect 740 15573 840 15673
rect 740 15373 840 15473
rect 740 15173 840 15273
rect 740 14973 840 15073
rect 1235 17373 1335 17473
rect 1235 17173 1335 17273
rect 1235 16973 1335 17073
rect 1235 16773 1335 16873
rect 1235 16573 1335 16673
rect 1235 16373 1335 16473
rect 1235 16173 1335 16273
rect 1235 15973 1335 16073
rect 1235 15773 1335 15873
rect 1235 15573 1335 15673
rect 1235 15373 1335 15473
rect 1235 15173 1335 15273
rect 1235 14973 1335 15073
rect 1740 17373 1840 17473
rect 1740 17173 1840 17273
rect 1740 16973 1840 17073
rect 1740 16773 1840 16873
rect 1740 16573 1840 16673
rect 1740 16373 1840 16473
rect 1740 16173 1840 16273
rect 1740 15973 1840 16073
rect 1740 15773 1840 15873
rect 1740 15573 1840 15673
rect 1740 15373 1840 15473
rect 1740 15173 1840 15273
rect 1740 14973 1840 15073
rect 2235 17373 2335 17473
rect 2235 17173 2335 17273
rect 2235 16973 2335 17073
rect 2235 16773 2335 16873
rect 2235 16573 2335 16673
rect 2235 16373 2335 16473
rect 2235 16173 2335 16273
rect 2235 15973 2335 16073
rect 2235 15773 2335 15873
rect 2235 15573 2335 15673
rect 2235 15373 2335 15473
rect 2235 15173 2335 15273
rect 2235 14973 2335 15073
rect 2740 17373 2840 17473
rect 2740 17173 2840 17273
rect 2740 16973 2840 17073
rect 2740 16773 2840 16873
rect 2740 16573 2840 16673
rect 2740 16373 2840 16473
rect 2740 16173 2840 16273
rect 2740 15973 2840 16073
rect 2740 15773 2840 15873
rect 2740 15573 2840 15673
rect 2740 15373 2840 15473
rect 2740 15173 2840 15273
rect 2740 14973 2840 15073
rect 3235 17373 3335 17473
rect 3235 17173 3335 17273
rect 3235 16973 3335 17073
rect 3235 16773 3335 16873
rect 3235 16573 3335 16673
rect 3235 16373 3335 16473
rect 3235 16173 3335 16273
rect 3235 15973 3335 16073
rect 3235 15773 3335 15873
rect 3235 15573 3335 15673
rect 3235 15373 3335 15473
rect 3235 15173 3335 15273
rect 3235 14973 3335 15073
rect 3740 17373 3840 17473
rect 3740 17173 3840 17273
rect 3740 16973 3840 17073
rect 3740 16773 3840 16873
rect 3740 16573 3840 16673
rect 3740 16373 3840 16473
rect 3740 16173 3840 16273
rect 3740 15973 3840 16073
rect 3740 15773 3840 15873
rect 3740 15573 3840 15673
rect 3740 15373 3840 15473
rect 3740 15173 3840 15273
rect 3740 14973 3840 15073
rect 4235 17373 4335 17473
rect 4235 17173 4335 17273
rect 4235 16973 4335 17073
rect 4235 16773 4335 16873
rect 4235 16573 4335 16673
rect 4235 16373 4335 16473
rect 4235 16173 4335 16273
rect 4235 15973 4335 16073
rect 4235 15773 4335 15873
rect 4235 15573 4335 15673
rect 4235 15373 4335 15473
rect 4235 15173 4335 15273
rect 4235 14973 4335 15073
rect 4740 17373 4840 17473
rect 4740 17173 4840 17273
rect 4740 16973 4840 17073
rect 4740 16773 4840 16873
rect 4740 16573 4840 16673
rect 4740 16373 4840 16473
rect 4740 16173 4840 16273
rect 4740 15973 4840 16073
rect 4740 15773 4840 15873
rect 4740 15573 4840 15673
rect 4740 15373 4840 15473
rect 4740 15173 4840 15273
rect 4740 14973 4840 15073
rect 5235 17373 5335 17473
rect 5235 17173 5335 17273
rect 5235 16973 5335 17073
rect 5235 16773 5335 16873
rect 5235 16573 5335 16673
rect 5235 16373 5335 16473
rect 5235 16173 5335 16273
rect 5235 15973 5335 16073
rect 5235 15773 5335 15873
rect 5235 15573 5335 15673
rect 5235 15373 5335 15473
rect 5235 15173 5335 15273
rect 5235 14973 5335 15073
rect 5740 17373 5840 17473
rect 5740 17173 5840 17273
rect 5740 16973 5840 17073
rect 5740 16773 5840 16873
rect 5740 16573 5840 16673
rect 5740 16373 5840 16473
rect 5740 16173 5840 16273
rect 5740 15973 5840 16073
rect 5740 15773 5840 15873
rect 5740 15573 5840 15673
rect 5740 15373 5840 15473
rect 5740 15173 5840 15273
rect 5740 14973 5840 15073
rect 6235 17373 6335 17473
rect 6235 17173 6335 17273
rect 6235 16973 6335 17073
rect 6235 16773 6335 16873
rect 6235 16573 6335 16673
rect 6235 16373 6335 16473
rect 6235 16173 6335 16273
rect 6235 15973 6335 16073
rect 6235 15773 6335 15873
rect 6235 15573 6335 15673
rect 6235 15373 6335 15473
rect 6235 15173 6335 15273
rect 6235 14973 6335 15073
rect 6740 17373 6840 17473
rect 6740 17173 6840 17273
rect 6740 16973 6840 17073
rect 6740 16773 6840 16873
rect 6740 16573 6840 16673
rect 6740 16373 6840 16473
rect 6740 16173 6840 16273
rect 6740 15973 6840 16073
rect 6740 15773 6840 15873
rect 6740 15573 6840 15673
rect 6740 15373 6840 15473
rect 6740 15173 6840 15273
rect 6740 14973 6840 15073
rect 7235 17373 7335 17473
rect 7235 17173 7335 17273
rect 7235 16973 7335 17073
rect 7235 16773 7335 16873
rect 7235 16573 7335 16673
rect 7235 16373 7335 16473
rect 7235 16173 7335 16273
rect 7235 15973 7335 16073
rect 7235 15773 7335 15873
rect 7235 15573 7335 15673
rect 7235 15373 7335 15473
rect 7235 15173 7335 15273
rect 7235 14973 7335 15073
rect 7740 17373 7840 17473
rect 7740 17173 7840 17273
rect 7740 16973 7840 17073
rect 7740 16773 7840 16873
rect 7740 16573 7840 16673
rect 7740 16373 7840 16473
rect 7740 16173 7840 16273
rect 7740 15973 7840 16073
rect 7740 15773 7840 15873
rect 7740 15573 7840 15673
rect 7740 15373 7840 15473
rect 7740 15173 7840 15273
rect 7740 14973 7840 15073
rect 8235 17373 8335 17473
rect 8235 17173 8335 17273
rect 8235 16973 8335 17073
rect 8235 16773 8335 16873
rect 8235 16573 8335 16673
rect 8235 16373 8335 16473
rect 8235 16173 8335 16273
rect 8235 15973 8335 16073
rect 8235 15773 8335 15873
rect 8235 15573 8335 15673
rect 8235 15373 8335 15473
rect 8235 15173 8335 15273
rect 8235 14973 8335 15073
rect 8740 17373 8840 17473
rect 8740 17173 8840 17273
rect 8740 16973 8840 17073
rect 8740 16773 8840 16873
rect 8740 16573 8840 16673
rect 8740 16373 8840 16473
rect 8740 16173 8840 16273
rect 8740 15973 8840 16073
rect 8740 15773 8840 15873
rect 8740 15573 8840 15673
rect 8740 15373 8840 15473
rect 8740 15173 8840 15273
rect 8740 14973 8840 15073
rect 9235 17373 9335 17473
rect 9235 17173 9335 17273
rect 9235 16973 9335 17073
rect 9235 16773 9335 16873
rect 9235 16573 9335 16673
rect 9235 16373 9335 16473
rect 9235 16173 9335 16273
rect 9235 15973 9335 16073
rect 9235 15773 9335 15873
rect 9235 15573 9335 15673
rect 9235 15373 9335 15473
rect 9235 15173 9335 15273
rect 9235 14973 9335 15073
rect 9740 17373 9840 17473
rect 9740 17173 9840 17273
rect 9740 16973 9840 17073
rect 9740 16773 9840 16873
rect 9740 16573 9840 16673
rect 9740 16373 9840 16473
rect 9740 16173 9840 16273
rect 9740 15973 9840 16073
rect 9740 15773 9840 15873
rect 9740 15573 9840 15673
rect 9740 15373 9840 15473
rect 9740 15173 9840 15273
rect 9740 14973 9840 15073
rect -242 11646 -142 11746
rect -242 11446 -142 11546
rect -242 11246 -142 11346
rect -242 11046 -142 11146
rect -242 10846 -142 10946
rect -242 10646 -142 10746
rect -242 10446 -142 10546
rect -242 10246 -142 10346
rect -242 10046 -142 10146
rect -242 9846 -142 9946
rect -242 9646 -142 9746
rect -242 9446 -142 9546
rect -242 9246 -142 9346
rect 263 11646 363 11746
rect 263 11446 363 11546
rect 263 11246 363 11346
rect 263 11046 363 11146
rect 263 10846 363 10946
rect 263 10646 363 10746
rect 263 10446 363 10546
rect 263 10246 363 10346
rect 263 10046 363 10146
rect 263 9846 363 9946
rect 263 9646 363 9746
rect 263 9446 363 9546
rect 263 9246 363 9346
rect 758 11646 858 11746
rect 758 11446 858 11546
rect 758 11246 858 11346
rect 758 11046 858 11146
rect 758 10846 858 10946
rect 758 10646 858 10746
rect 758 10446 858 10546
rect 758 10246 858 10346
rect 758 10046 858 10146
rect 758 9846 858 9946
rect 758 9646 858 9746
rect 758 9446 858 9546
rect 758 9246 858 9346
rect 1263 11646 1363 11746
rect 1263 11446 1363 11546
rect 1263 11246 1363 11346
rect 1263 11046 1363 11146
rect 1263 10846 1363 10946
rect 1263 10646 1363 10746
rect 1263 10446 1363 10546
rect 1263 10246 1363 10346
rect 1263 10046 1363 10146
rect 1263 9846 1363 9946
rect 1263 9646 1363 9746
rect 1263 9446 1363 9546
rect 1263 9246 1363 9346
rect 1758 11646 1858 11746
rect 1758 11446 1858 11546
rect 1758 11246 1858 11346
rect 1758 11046 1858 11146
rect 1758 10846 1858 10946
rect 1758 10646 1858 10746
rect 1758 10446 1858 10546
rect 1758 10246 1858 10346
rect 1758 10046 1858 10146
rect 1758 9846 1858 9946
rect 1758 9646 1858 9746
rect 1758 9446 1858 9546
rect 1758 9246 1858 9346
rect 2263 11646 2363 11746
rect 2263 11446 2363 11546
rect 2263 11246 2363 11346
rect 2263 11046 2363 11146
rect 2263 10846 2363 10946
rect 2263 10646 2363 10746
rect 2263 10446 2363 10546
rect 2263 10246 2363 10346
rect 2263 10046 2363 10146
rect 2263 9846 2363 9946
rect 2263 9646 2363 9746
rect 2263 9446 2363 9546
rect 2263 9246 2363 9346
rect 2758 11646 2858 11746
rect 2758 11446 2858 11546
rect 2758 11246 2858 11346
rect 2758 11046 2858 11146
rect 2758 10846 2858 10946
rect 2758 10646 2858 10746
rect 2758 10446 2858 10546
rect 2758 10246 2858 10346
rect 2758 10046 2858 10146
rect 2758 9846 2858 9946
rect 2758 9646 2858 9746
rect 2758 9446 2858 9546
rect 2758 9246 2858 9346
rect 3263 11646 3363 11746
rect 3263 11446 3363 11546
rect 3263 11246 3363 11346
rect 3263 11046 3363 11146
rect 3263 10846 3363 10946
rect 3263 10646 3363 10746
rect 3263 10446 3363 10546
rect 3263 10246 3363 10346
rect 3263 10046 3363 10146
rect 3263 9846 3363 9946
rect 3263 9646 3363 9746
rect 3263 9446 3363 9546
rect 3263 9246 3363 9346
rect 3758 11646 3858 11746
rect 3758 11446 3858 11546
rect 3758 11246 3858 11346
rect 3758 11046 3858 11146
rect 3758 10846 3858 10946
rect 3758 10646 3858 10746
rect 3758 10446 3858 10546
rect 3758 10246 3858 10346
rect 3758 10046 3858 10146
rect 3758 9846 3858 9946
rect 3758 9646 3858 9746
rect 3758 9446 3858 9546
rect 3758 9246 3858 9346
rect 4263 11646 4363 11746
rect 4263 11446 4363 11546
rect 4263 11246 4363 11346
rect 4263 11046 4363 11146
rect 4263 10846 4363 10946
rect 4263 10646 4363 10746
rect 4263 10446 4363 10546
rect 4263 10246 4363 10346
rect 4263 10046 4363 10146
rect 4263 9846 4363 9946
rect 4263 9646 4363 9746
rect 4263 9446 4363 9546
rect 4263 9246 4363 9346
rect 4758 11646 4858 11746
rect 4758 11446 4858 11546
rect 4758 11246 4858 11346
rect 4758 11046 4858 11146
rect 4758 10846 4858 10946
rect 4758 10646 4858 10746
rect 4758 10446 4858 10546
rect 4758 10246 4858 10346
rect 4758 10046 4858 10146
rect 4758 9846 4858 9946
rect 4758 9646 4858 9746
rect 4758 9446 4858 9546
rect 4758 9246 4858 9346
rect 5263 11646 5363 11746
rect 5263 11446 5363 11546
rect 5263 11246 5363 11346
rect 5263 11046 5363 11146
rect 5263 10846 5363 10946
rect 5263 10646 5363 10746
rect 5263 10446 5363 10546
rect 5263 10246 5363 10346
rect 5263 10046 5363 10146
rect 5263 9846 5363 9946
rect 5263 9646 5363 9746
rect 5263 9446 5363 9546
rect 5263 9246 5363 9346
rect 5758 11646 5858 11746
rect 5758 11446 5858 11546
rect 5758 11246 5858 11346
rect 5758 11046 5858 11146
rect 5758 10846 5858 10946
rect 5758 10646 5858 10746
rect 5758 10446 5858 10546
rect 5758 10246 5858 10346
rect 5758 10046 5858 10146
rect 5758 9846 5858 9946
rect 5758 9646 5858 9746
rect 5758 9446 5858 9546
rect 5758 9246 5858 9346
rect 6263 11646 6363 11746
rect 6263 11446 6363 11546
rect 6263 11246 6363 11346
rect 6263 11046 6363 11146
rect 6263 10846 6363 10946
rect 6263 10646 6363 10746
rect 6263 10446 6363 10546
rect 6263 10246 6363 10346
rect 6263 10046 6363 10146
rect 6263 9846 6363 9946
rect 6263 9646 6363 9746
rect 6263 9446 6363 9546
rect 6263 9246 6363 9346
rect 6758 11646 6858 11746
rect 6758 11446 6858 11546
rect 6758 11246 6858 11346
rect 6758 11046 6858 11146
rect 6758 10846 6858 10946
rect 6758 10646 6858 10746
rect 6758 10446 6858 10546
rect 6758 10246 6858 10346
rect 6758 10046 6858 10146
rect 6758 9846 6858 9946
rect 6758 9646 6858 9746
rect 6758 9446 6858 9546
rect 6758 9246 6858 9346
rect 7263 11646 7363 11746
rect 7263 11446 7363 11546
rect 7263 11246 7363 11346
rect 7263 11046 7363 11146
rect 7263 10846 7363 10946
rect 7263 10646 7363 10746
rect 7263 10446 7363 10546
rect 7263 10246 7363 10346
rect 7263 10046 7363 10146
rect 7263 9846 7363 9946
rect 7263 9646 7363 9746
rect 7263 9446 7363 9546
rect 7263 9246 7363 9346
rect 7758 11646 7858 11746
rect 7758 11446 7858 11546
rect 7758 11246 7858 11346
rect 7758 11046 7858 11146
rect 7758 10846 7858 10946
rect 7758 10646 7858 10746
rect 7758 10446 7858 10546
rect 7758 10246 7858 10346
rect 7758 10046 7858 10146
rect 7758 9846 7858 9946
rect 7758 9646 7858 9746
rect 7758 9446 7858 9546
rect 7758 9246 7858 9346
rect 8263 11646 8363 11746
rect 8263 11446 8363 11546
rect 8263 11246 8363 11346
rect 8263 11046 8363 11146
rect 8263 10846 8363 10946
rect 8263 10646 8363 10746
rect 8263 10446 8363 10546
rect 8263 10246 8363 10346
rect 8263 10046 8363 10146
rect 8263 9846 8363 9946
rect 8263 9646 8363 9746
rect 8263 9446 8363 9546
rect 8263 9246 8363 9346
rect 8758 11646 8858 11746
rect 8758 11446 8858 11546
rect 8758 11246 8858 11346
rect 8758 11046 8858 11146
rect 8758 10846 8858 10946
rect 8758 10646 8858 10746
rect 8758 10446 8858 10546
rect 8758 10246 8858 10346
rect 8758 10046 8858 10146
rect 8758 9846 8858 9946
rect 8758 9646 8858 9746
rect 8758 9446 8858 9546
rect 8758 9246 8858 9346
rect 9263 11646 9363 11746
rect 9263 11446 9363 11546
rect 9263 11246 9363 11346
rect 9263 11046 9363 11146
rect 9263 10846 9363 10946
rect 9263 10646 9363 10746
rect 9263 10446 9363 10546
rect 9263 10246 9363 10346
rect 9263 10046 9363 10146
rect 9263 9846 9363 9946
rect 9263 9646 9363 9746
rect 9263 9446 9363 9546
rect 9263 9246 9363 9346
rect 9782 11642 9882 11742
rect 9782 11442 9882 11542
rect 9782 11242 9882 11342
rect 9782 11042 9882 11142
rect 9782 10842 9882 10942
rect 9782 10642 9882 10742
rect 9782 10442 9882 10542
rect 9782 10242 9882 10342
rect 9782 10042 9882 10142
rect 9782 9842 9882 9942
rect 9782 9642 9882 9742
rect 9782 9442 9882 9542
rect 9782 9242 9882 9342
<< psubdiff >>
rect 2259 6743 2524 6796
rect 2259 6555 2313 6743
rect 2481 6555 2524 6743
rect 2259 6496 2524 6555
<< nsubdiff >>
rect 9801 14330 10208 14367
rect 9801 14144 9851 14330
rect 10161 14144 10208 14330
rect 9801 14097 10208 14144
rect 9865 12599 10221 12650
rect 9865 12401 9911 12599
rect 10175 12401 10221 12599
rect 9865 12342 10221 12401
<< psubdiffcont >>
rect 2313 6555 2481 6743
<< nsubdiffcont >>
rect 9851 14144 10161 14330
rect 9911 12401 10175 12599
<< poly >>
rect -11 18166 89 18186
rect -11 18079 0 18166
rect 76 18079 89 18166
rect -11 17707 89 18079
rect 489 18166 589 18186
rect 489 18079 500 18166
rect 576 18079 589 18166
rect 489 17707 589 18079
rect 989 18166 1089 18186
rect 989 18079 1000 18166
rect 1076 18079 1089 18166
rect 989 17707 1089 18079
rect 1489 18166 1589 18186
rect 1489 18079 1500 18166
rect 1576 18079 1589 18166
rect 1489 17707 1589 18079
rect 1989 18166 2089 18186
rect 1989 18079 2000 18166
rect 2076 18079 2089 18166
rect 1989 17707 2089 18079
rect 2489 18166 2589 18186
rect 2489 18079 2500 18166
rect 2576 18079 2589 18166
rect 2489 17707 2589 18079
rect 2989 18166 3089 18186
rect 2989 18079 3000 18166
rect 3076 18079 3089 18166
rect 2989 17707 3089 18079
rect 3489 18166 3589 18186
rect 3489 18079 3500 18166
rect 3576 18079 3589 18166
rect 3489 17707 3589 18079
rect 3989 18166 4089 18186
rect 3989 18079 4000 18166
rect 4076 18079 4089 18166
rect 3989 17707 4089 18079
rect 4489 18166 4589 18186
rect 4489 18079 4500 18166
rect 4576 18079 4589 18166
rect 4489 17707 4589 18079
rect 4989 18166 5089 18186
rect 4989 18079 5000 18166
rect 5076 18079 5089 18166
rect 4989 17707 5089 18079
rect 5489 18166 5589 18186
rect 5489 18079 5500 18166
rect 5576 18079 5589 18166
rect 5489 17707 5589 18079
rect 5989 18166 6089 18186
rect 5989 18079 6000 18166
rect 6076 18079 6089 18166
rect 5989 17707 6089 18079
rect 6489 18166 6589 18186
rect 6489 18079 6500 18166
rect 6576 18079 6589 18166
rect 6489 17707 6589 18079
rect 6989 18166 7089 18186
rect 6989 18079 7000 18166
rect 7076 18079 7089 18166
rect 6989 17707 7089 18079
rect 7489 18166 7589 18186
rect 7489 18079 7500 18166
rect 7576 18079 7589 18166
rect 7489 17707 7589 18079
rect 7989 18166 8089 18186
rect 7989 18079 8000 18166
rect 8076 18079 8089 18166
rect 7989 17707 8089 18079
rect 8489 18166 8589 18186
rect 8489 18079 8500 18166
rect 8576 18079 8589 18166
rect 8489 17707 8589 18079
rect 8989 18166 9089 18186
rect 8989 18079 9000 18166
rect 9076 18079 9089 18166
rect 8989 17707 9089 18079
rect 9489 18166 9589 18186
rect 9489 18079 9500 18166
rect 9576 18079 9589 18166
rect 9489 17707 9589 18079
rect -11 14317 89 14707
rect -1235 14302 89 14317
rect -1249 14291 89 14302
rect 489 14291 589 14707
rect 989 14291 1089 14707
rect 1489 14291 1589 14707
rect 1989 14291 2089 14707
rect 2489 14291 2589 14707
rect 2989 14291 3089 14707
rect 3489 14291 3589 14707
rect 3989 14291 4089 14707
rect 4489 14291 4589 14707
rect 4989 14291 5089 14707
rect 5489 14291 5589 14707
rect 5989 14291 6089 14707
rect 6489 14291 6589 14707
rect 6989 14291 7089 14707
rect 7489 14291 7589 14707
rect 7989 14291 8089 14707
rect 8489 14291 8589 14707
rect 8989 14291 9089 14707
rect 9489 14291 9589 14707
rect -1249 14100 9589 14291
rect -1249 13878 -730 14100
rect -11 14091 9589 14100
rect -1249 13178 -1214 13878
rect -765 13178 -730 13878
rect -1249 13092 -730 13178
rect 5034 12628 5448 14091
rect 9 12428 9609 12628
rect 9 12012 109 12428
rect 509 12012 609 12428
rect 1009 12012 1109 12428
rect 1509 12012 1609 12428
rect 2009 12012 2109 12428
rect 2509 12012 2609 12428
rect 3009 12012 3109 12428
rect 3509 12012 3609 12428
rect 4009 12012 4109 12428
rect 4509 12012 4609 12428
rect 5009 12423 5448 12428
rect 5009 12012 5109 12423
rect 5509 12012 5609 12428
rect 6009 12012 6109 12428
rect 6509 12012 6609 12428
rect 7009 12012 7109 12428
rect 7509 12012 7609 12428
rect 8009 12012 8109 12428
rect 8509 12012 8609 12428
rect 9009 12012 9109 12428
rect 9509 12012 9609 12428
rect 9 8533 109 9012
rect 509 8533 609 9012
rect 1009 8533 1109 9012
rect 1509 8533 1609 9012
rect 2009 8533 2109 9012
rect 2509 8533 2609 9012
rect 3009 8533 3109 9012
rect 3509 8533 3609 9012
rect 4009 8533 4109 9012
rect 4509 8533 4609 9012
rect 5009 8533 5109 9012
rect 5509 8533 5609 9012
rect 6009 8533 6109 9012
rect 6509 8533 6609 9012
rect 7009 8533 7109 9012
rect 7509 8533 7609 9012
rect 8009 8533 8109 9012
rect 8509 8533 8609 9012
rect 9009 8533 9109 9012
rect 9509 8533 9609 9012
rect -146 7343 149 7373
rect -146 7101 -124 7343
rect 118 7101 149 7343
rect -146 7073 149 7101
rect 49 7044 149 7073
rect 449 7044 549 7107
rect 849 7044 949 7107
rect 1249 7044 1349 7107
rect 1649 7044 1749 7107
rect 49 5807 149 5851
rect 449 5807 549 5851
rect 849 5807 949 5851
rect 1249 5807 1349 5851
rect 1649 5807 1749 5851
rect 49 5707 1749 5807
<< polycont >>
rect 0 18079 76 18166
rect 500 18079 576 18166
rect 1000 18079 1076 18166
rect 1500 18079 1576 18166
rect 2000 18079 2076 18166
rect 2500 18079 2576 18166
rect 3000 18079 3076 18166
rect 3500 18079 3576 18166
rect 4000 18079 4076 18166
rect 4500 18079 4576 18166
rect 5000 18079 5076 18166
rect 5500 18079 5576 18166
rect 6000 18079 6076 18166
rect 6500 18079 6576 18166
rect 7000 18079 7076 18166
rect 7500 18079 7576 18166
rect 8000 18079 8076 18166
rect 8500 18079 8576 18166
rect 9000 18079 9076 18166
rect 9500 18079 9576 18166
rect -1214 13178 -765 13878
rect -124 7101 118 7343
<< locali >>
rect 235 18186 335 18187
rect 1235 18186 1335 18187
rect 2235 18186 2335 18187
rect 3235 18186 3335 18187
rect 4235 18186 4335 18187
rect 5235 18186 5335 18187
rect 6235 18186 6335 18187
rect 7235 18186 7335 18187
rect 8235 18186 8335 18187
rect 9235 18186 9335 18187
rect -11 18166 9589 18186
rect -11 18079 0 18166
rect 76 18079 500 18166
rect 576 18079 1000 18166
rect 1076 18079 1500 18166
rect 1576 18079 2000 18166
rect 2076 18079 2500 18166
rect 2576 18079 3000 18166
rect 3076 18079 3500 18166
rect 3576 18079 4000 18166
rect 4076 18079 4500 18166
rect 4576 18079 5000 18166
rect 5076 18079 5500 18166
rect 5576 18079 6000 18166
rect 6076 18079 6500 18166
rect 6576 18079 7000 18166
rect 7076 18079 7500 18166
rect 7576 18079 8000 18166
rect 8076 18079 8500 18166
rect 8576 18079 9000 18166
rect 9076 18079 9500 18166
rect 9576 18079 9589 18166
rect -11 18055 9589 18079
rect -284 17477 -184 17557
rect -284 17277 -184 17377
rect -284 17077 -184 17177
rect -284 16877 -184 16977
rect -284 16677 -184 16777
rect -284 16477 -184 16577
rect -284 16277 -184 16377
rect -284 16077 -184 16177
rect -284 15877 -184 15977
rect -284 15677 -184 15777
rect -284 15477 -184 15577
rect -284 15277 -184 15377
rect -284 15077 -184 15177
rect -1249 13878 -730 14001
rect -1249 13178 -1214 13878
rect -765 13178 -730 13878
rect -284 13760 -184 14977
rect 235 17473 335 18055
rect 235 17273 335 17373
rect 235 17073 335 17173
rect 235 16873 335 16973
rect 235 16673 335 16773
rect 235 16473 335 16573
rect 235 16273 335 16373
rect 235 16073 335 16173
rect 235 15873 335 15973
rect 235 15673 335 15773
rect 235 15473 335 15573
rect 235 15273 335 15373
rect 235 15073 335 15173
rect 235 14813 335 14973
rect 740 17473 840 17514
rect 740 17273 840 17373
rect 740 17073 840 17173
rect 740 16873 840 16973
rect 740 16673 840 16773
rect 740 16473 840 16573
rect 740 16273 840 16373
rect 740 16073 840 16173
rect 740 15873 840 15973
rect 740 15673 840 15773
rect 740 15473 840 15573
rect 740 15273 840 15373
rect 740 15073 840 15173
rect 740 13760 840 14973
rect 1235 17473 1335 18055
rect 1235 17273 1335 17373
rect 1235 17073 1335 17173
rect 1235 16873 1335 16973
rect 1235 16673 1335 16773
rect 1235 16473 1335 16573
rect 1235 16273 1335 16373
rect 1235 16073 1335 16173
rect 1235 15873 1335 15973
rect 1235 15673 1335 15773
rect 1235 15473 1335 15573
rect 1235 15273 1335 15373
rect 1235 15073 1335 15173
rect 1235 14813 1335 14973
rect 1740 17473 1840 17514
rect 1740 17273 1840 17373
rect 1740 17073 1840 17173
rect 1740 16873 1840 16973
rect 1740 16673 1840 16773
rect 1740 16473 1840 16573
rect 1740 16273 1840 16373
rect 1740 16073 1840 16173
rect 1740 15873 1840 15973
rect 1740 15673 1840 15773
rect 1740 15473 1840 15573
rect 1740 15273 1840 15373
rect 1740 15073 1840 15173
rect 1740 13760 1840 14973
rect 2235 17473 2335 18055
rect 2235 17273 2335 17373
rect 2235 17073 2335 17173
rect 2235 16873 2335 16973
rect 2235 16673 2335 16773
rect 2235 16473 2335 16573
rect 2235 16273 2335 16373
rect 2235 16073 2335 16173
rect 2235 15873 2335 15973
rect 2235 15673 2335 15773
rect 2235 15473 2335 15573
rect 2235 15273 2335 15373
rect 2235 15073 2335 15173
rect 2235 14813 2335 14973
rect 2740 17473 2840 17514
rect 2740 17273 2840 17373
rect 2740 17073 2840 17173
rect 2740 16873 2840 16973
rect 2740 16673 2840 16773
rect 2740 16473 2840 16573
rect 2740 16273 2840 16373
rect 2740 16073 2840 16173
rect 2740 15873 2840 15973
rect 2740 15673 2840 15773
rect 2740 15473 2840 15573
rect 2740 15273 2840 15373
rect 2740 15073 2840 15173
rect 2740 13760 2840 14973
rect 3235 17473 3335 18055
rect 3235 17273 3335 17373
rect 3235 17073 3335 17173
rect 3235 16873 3335 16973
rect 3235 16673 3335 16773
rect 3235 16473 3335 16573
rect 3235 16273 3335 16373
rect 3235 16073 3335 16173
rect 3235 15873 3335 15973
rect 3235 15673 3335 15773
rect 3235 15473 3335 15573
rect 3235 15273 3335 15373
rect 3235 15073 3335 15173
rect 3235 14813 3335 14973
rect 3740 17473 3840 17514
rect 3740 17273 3840 17373
rect 3740 17073 3840 17173
rect 3740 16873 3840 16973
rect 3740 16673 3840 16773
rect 3740 16473 3840 16573
rect 3740 16273 3840 16373
rect 3740 16073 3840 16173
rect 3740 15873 3840 15973
rect 3740 15673 3840 15773
rect 3740 15473 3840 15573
rect 3740 15273 3840 15373
rect 3740 15073 3840 15173
rect 3740 13760 3840 14973
rect 4235 17473 4335 18055
rect 4235 17273 4335 17373
rect 4235 17073 4335 17173
rect 4235 16873 4335 16973
rect 4235 16673 4335 16773
rect 4235 16473 4335 16573
rect 4235 16273 4335 16373
rect 4235 16073 4335 16173
rect 4235 15873 4335 15973
rect 4235 15673 4335 15773
rect 4235 15473 4335 15573
rect 4235 15273 4335 15373
rect 4235 15073 4335 15173
rect 4235 14813 4335 14973
rect 4740 17473 4840 17514
rect 4740 17273 4840 17373
rect 4740 17073 4840 17173
rect 4740 16873 4840 16973
rect 4740 16673 4840 16773
rect 4740 16473 4840 16573
rect 4740 16273 4840 16373
rect 4740 16073 4840 16173
rect 4740 15873 4840 15973
rect 4740 15673 4840 15773
rect 4740 15473 4840 15573
rect 4740 15273 4840 15373
rect 4740 15073 4840 15173
rect 4740 13760 4840 14973
rect 5235 17473 5335 18055
rect 5235 17273 5335 17373
rect 5235 17073 5335 17173
rect 5235 16873 5335 16973
rect 5235 16673 5335 16773
rect 5235 16473 5335 16573
rect 5235 16273 5335 16373
rect 5235 16073 5335 16173
rect 5235 15873 5335 15973
rect 5235 15673 5335 15773
rect 5235 15473 5335 15573
rect 5235 15273 5335 15373
rect 5235 15073 5335 15173
rect 5235 14813 5335 14973
rect 5740 17473 5840 17514
rect 5740 17273 5840 17373
rect 5740 17073 5840 17173
rect 5740 16873 5840 16973
rect 5740 16673 5840 16773
rect 5740 16473 5840 16573
rect 5740 16273 5840 16373
rect 5740 16073 5840 16173
rect 5740 15873 5840 15973
rect 5740 15673 5840 15773
rect 5740 15473 5840 15573
rect 5740 15273 5840 15373
rect 5740 15073 5840 15173
rect 5740 13760 5840 14973
rect 6235 17473 6335 18055
rect 6235 17273 6335 17373
rect 6235 17073 6335 17173
rect 6235 16873 6335 16973
rect 6235 16673 6335 16773
rect 6235 16473 6335 16573
rect 6235 16273 6335 16373
rect 6235 16073 6335 16173
rect 6235 15873 6335 15973
rect 6235 15673 6335 15773
rect 6235 15473 6335 15573
rect 6235 15273 6335 15373
rect 6235 15073 6335 15173
rect 6235 14813 6335 14973
rect 6740 17473 6840 17514
rect 6740 17273 6840 17373
rect 6740 17073 6840 17173
rect 6740 16873 6840 16973
rect 6740 16673 6840 16773
rect 6740 16473 6840 16573
rect 6740 16273 6840 16373
rect 6740 16073 6840 16173
rect 6740 15873 6840 15973
rect 6740 15673 6840 15773
rect 6740 15473 6840 15573
rect 6740 15273 6840 15373
rect 6740 15073 6840 15173
rect 6740 13760 6840 14973
rect 7235 17473 7335 18055
rect 7235 17273 7335 17373
rect 7235 17073 7335 17173
rect 7235 16873 7335 16973
rect 7235 16673 7335 16773
rect 7235 16473 7335 16573
rect 7235 16273 7335 16373
rect 7235 16073 7335 16173
rect 7235 15873 7335 15973
rect 7235 15673 7335 15773
rect 7235 15473 7335 15573
rect 7235 15273 7335 15373
rect 7235 15073 7335 15173
rect 7235 14813 7335 14973
rect 7740 17473 7840 17514
rect 7740 17273 7840 17373
rect 7740 17073 7840 17173
rect 7740 16873 7840 16973
rect 7740 16673 7840 16773
rect 7740 16473 7840 16573
rect 7740 16273 7840 16373
rect 7740 16073 7840 16173
rect 7740 15873 7840 15973
rect 7740 15673 7840 15773
rect 7740 15473 7840 15573
rect 7740 15273 7840 15373
rect 7740 15073 7840 15173
rect 7740 13760 7840 14973
rect 8235 17473 8335 18055
rect 8235 17273 8335 17373
rect 8235 17073 8335 17173
rect 8235 16873 8335 16973
rect 8235 16673 8335 16773
rect 8235 16473 8335 16573
rect 8235 16273 8335 16373
rect 8235 16073 8335 16173
rect 8235 15873 8335 15973
rect 8235 15673 8335 15773
rect 8235 15473 8335 15573
rect 8235 15273 8335 15373
rect 8235 15073 8335 15173
rect 8235 14813 8335 14973
rect 8740 17473 8840 17514
rect 8740 17273 8840 17373
rect 8740 17073 8840 17173
rect 8740 16873 8840 16973
rect 8740 16673 8840 16773
rect 8740 16473 8840 16573
rect 8740 16273 8840 16373
rect 8740 16073 8840 16173
rect 8740 15873 8840 15973
rect 8740 15673 8840 15773
rect 8740 15473 8840 15573
rect 8740 15273 8840 15373
rect 8740 15073 8840 15173
rect 8740 13760 8840 14973
rect 9235 17473 9335 18055
rect 9235 17273 9335 17373
rect 9235 17073 9335 17173
rect 9235 16873 9335 16973
rect 9235 16673 9335 16773
rect 9235 16473 9335 16573
rect 9235 16273 9335 16373
rect 9235 16073 9335 16173
rect 9235 15873 9335 15973
rect 9235 15673 9335 15773
rect 9235 15473 9335 15573
rect 9235 15273 9335 15373
rect 9235 15073 9335 15173
rect 9235 14813 9335 14973
rect 9740 17473 9840 17514
rect 9740 17273 9840 17373
rect 9740 17073 9840 17173
rect 9740 16873 9840 16973
rect 9740 16673 9840 16773
rect 9740 16473 9840 16573
rect 9740 16273 9840 16373
rect 9740 16073 9840 16173
rect 9740 15873 9840 15973
rect 9740 15673 9840 15773
rect 9740 15473 9840 15573
rect 9740 15273 9840 15373
rect 9740 15073 9840 15173
rect -388 13738 8840 13760
rect 9740 14471 9840 14973
rect 9740 14330 10285 14471
rect 9740 14144 9851 14330
rect 10161 14144 10285 14330
rect 9740 13738 10285 14144
rect -388 13726 10285 13738
rect -388 13557 10577 13726
rect -388 13535 9933 13557
rect -236 13206 65 13535
rect 710 13513 9933 13535
rect -1249 13092 -730 13178
rect -242 13184 8888 13206
rect 9415 13184 9933 13513
rect -242 13171 9933 13184
rect 10404 13171 10577 13557
rect -242 12981 10577 13171
rect -242 11746 -142 12981
rect 758 12959 10577 12981
rect -242 11546 -142 11646
rect -242 11346 -142 11446
rect -242 11146 -142 11246
rect -242 10946 -142 11046
rect -242 10746 -142 10846
rect -242 10546 -142 10646
rect -242 10346 -142 10446
rect -242 10146 -142 10246
rect -242 9946 -142 10046
rect -242 9746 -142 9846
rect -242 9546 -142 9646
rect -242 9346 -142 9446
rect -242 9205 -142 9246
rect 263 11746 363 11906
rect 263 11546 363 11646
rect 263 11346 363 11446
rect 263 11146 363 11246
rect 263 10946 363 11046
rect 263 10746 363 10846
rect 263 10546 363 10646
rect 263 10346 363 10446
rect 263 10146 363 10246
rect 263 9946 363 10046
rect 263 9746 363 9846
rect 263 9546 363 9646
rect 263 9346 363 9446
rect 263 8130 363 9246
rect 758 11746 858 12959
rect 758 11546 858 11646
rect 758 11346 858 11446
rect 758 11146 858 11246
rect 758 10946 858 11046
rect 758 10746 858 10846
rect 758 10546 858 10646
rect 758 10346 858 10446
rect 758 10146 858 10246
rect 758 9946 858 10046
rect 758 9746 858 9846
rect 758 9546 858 9646
rect 758 9346 858 9446
rect 758 9205 858 9246
rect 1263 11746 1363 11906
rect 1263 11546 1363 11646
rect 1263 11346 1363 11446
rect 1263 11146 1363 11246
rect 1263 10946 1363 11046
rect 1263 10746 1363 10846
rect 1263 10546 1363 10646
rect 1263 10346 1363 10446
rect 1263 10146 1363 10246
rect 1263 9946 1363 10046
rect 1263 9746 1363 9846
rect 1263 9546 1363 9646
rect 1263 9346 1363 9446
rect 1263 8130 1363 9246
rect 1758 11746 1858 12959
rect 1758 11546 1858 11646
rect 1758 11346 1858 11446
rect 1758 11146 1858 11246
rect 1758 10946 1858 11046
rect 1758 10746 1858 10846
rect 1758 10546 1858 10646
rect 1758 10346 1858 10446
rect 1758 10146 1858 10246
rect 1758 9946 1858 10046
rect 1758 9746 1858 9846
rect 1758 9546 1858 9646
rect 1758 9346 1858 9446
rect 1758 9205 1858 9246
rect 2263 11746 2363 11906
rect 2263 11546 2363 11646
rect 2263 11346 2363 11446
rect 2263 11146 2363 11246
rect 2263 10946 2363 11046
rect 2263 10746 2363 10846
rect 2263 10546 2363 10646
rect 2263 10346 2363 10446
rect 2263 10146 2363 10246
rect 2263 9946 2363 10046
rect 2263 9746 2363 9846
rect 2263 9546 2363 9646
rect 2263 9346 2363 9446
rect 2263 8130 2363 9246
rect 2758 11746 2858 12959
rect 2758 11546 2858 11646
rect 2758 11346 2858 11446
rect 2758 11146 2858 11246
rect 2758 10946 2858 11046
rect 2758 10746 2858 10846
rect 2758 10546 2858 10646
rect 2758 10346 2858 10446
rect 2758 10146 2858 10246
rect 2758 9946 2858 10046
rect 2758 9746 2858 9846
rect 2758 9546 2858 9646
rect 2758 9346 2858 9446
rect 2758 9205 2858 9246
rect 3263 11746 3363 11906
rect 3263 11546 3363 11646
rect 3263 11346 3363 11446
rect 3263 11146 3363 11246
rect 3263 10946 3363 11046
rect 3263 10746 3363 10846
rect 3263 10546 3363 10646
rect 3263 10346 3363 10446
rect 3263 10146 3363 10246
rect 3263 9946 3363 10046
rect 3263 9746 3363 9846
rect 3263 9546 3363 9646
rect 3263 9346 3363 9446
rect 3263 8130 3363 9246
rect 3758 11746 3858 12959
rect 3758 11546 3858 11646
rect 3758 11346 3858 11446
rect 3758 11146 3858 11246
rect 3758 10946 3858 11046
rect 3758 10746 3858 10846
rect 3758 10546 3858 10646
rect 3758 10346 3858 10446
rect 3758 10146 3858 10246
rect 3758 9946 3858 10046
rect 3758 9746 3858 9846
rect 3758 9546 3858 9646
rect 3758 9346 3858 9446
rect 3758 9205 3858 9246
rect 4263 11746 4363 11906
rect 4263 11546 4363 11646
rect 4263 11346 4363 11446
rect 4263 11146 4363 11246
rect 4263 10946 4363 11046
rect 4263 10746 4363 10846
rect 4263 10546 4363 10646
rect 4263 10346 4363 10446
rect 4263 10146 4363 10246
rect 4263 9946 4363 10046
rect 4263 9746 4363 9846
rect 4263 9546 4363 9646
rect 4263 9346 4363 9446
rect 4263 8130 4363 9246
rect 4758 11746 4858 12959
rect 4758 11546 4858 11646
rect 4758 11346 4858 11446
rect 4758 11146 4858 11246
rect 4758 10946 4858 11046
rect 4758 10746 4858 10846
rect 4758 10546 4858 10646
rect 4758 10346 4858 10446
rect 4758 10146 4858 10246
rect 4758 9946 4858 10046
rect 4758 9746 4858 9846
rect 4758 9546 4858 9646
rect 4758 9346 4858 9446
rect 4758 9205 4858 9246
rect 5263 11746 5363 11906
rect 5263 11546 5363 11646
rect 5263 11346 5363 11446
rect 5263 11146 5363 11246
rect 5263 10946 5363 11046
rect 5263 10746 5363 10846
rect 5263 10546 5363 10646
rect 5263 10346 5363 10446
rect 5263 10146 5363 10246
rect 5263 9946 5363 10046
rect 5263 9746 5363 9846
rect 5263 9546 5363 9646
rect 5263 9346 5363 9446
rect 5263 8130 5363 9246
rect 5758 11746 5858 12959
rect 5758 11546 5858 11646
rect 5758 11346 5858 11446
rect 5758 11146 5858 11246
rect 5758 10946 5858 11046
rect 5758 10746 5858 10846
rect 5758 10546 5858 10646
rect 5758 10346 5858 10446
rect 5758 10146 5858 10246
rect 5758 9946 5858 10046
rect 5758 9746 5858 9846
rect 5758 9546 5858 9646
rect 5758 9346 5858 9446
rect 5758 9205 5858 9246
rect 6263 11746 6363 11906
rect 6263 11546 6363 11646
rect 6263 11346 6363 11446
rect 6263 11146 6363 11246
rect 6263 10946 6363 11046
rect 6263 10746 6363 10846
rect 6263 10546 6363 10646
rect 6263 10346 6363 10446
rect 6263 10146 6363 10246
rect 6263 9946 6363 10046
rect 6263 9746 6363 9846
rect 6263 9546 6363 9646
rect 6263 9346 6363 9446
rect 6263 8130 6363 9246
rect 6758 11746 6858 12959
rect 6758 11546 6858 11646
rect 6758 11346 6858 11446
rect 6758 11146 6858 11246
rect 6758 10946 6858 11046
rect 6758 10746 6858 10846
rect 6758 10546 6858 10646
rect 6758 10346 6858 10446
rect 6758 10146 6858 10246
rect 6758 9946 6858 10046
rect 6758 9746 6858 9846
rect 6758 9546 6858 9646
rect 6758 9346 6858 9446
rect 6758 9205 6858 9246
rect 7263 11746 7363 11906
rect 7263 11546 7363 11646
rect 7263 11346 7363 11446
rect 7263 11146 7363 11246
rect 7263 10946 7363 11046
rect 7263 10746 7363 10846
rect 7263 10546 7363 10646
rect 7263 10346 7363 10446
rect 7263 10146 7363 10246
rect 7263 9946 7363 10046
rect 7263 9746 7363 9846
rect 7263 9546 7363 9646
rect 7263 9346 7363 9446
rect 7263 8130 7363 9246
rect 7758 11746 7858 12959
rect 7758 11546 7858 11646
rect 7758 11346 7858 11446
rect 7758 11146 7858 11246
rect 7758 10946 7858 11046
rect 7758 10746 7858 10846
rect 7758 10546 7858 10646
rect 7758 10346 7858 10446
rect 7758 10146 7858 10246
rect 7758 9946 7858 10046
rect 7758 9746 7858 9846
rect 7758 9546 7858 9646
rect 7758 9346 7858 9446
rect 7758 9205 7858 9246
rect 8263 11746 8363 11906
rect 8263 11546 8363 11646
rect 8263 11346 8363 11446
rect 8263 11146 8363 11246
rect 8263 10946 8363 11046
rect 8263 10746 8363 10846
rect 8263 10546 8363 10646
rect 8263 10346 8363 10446
rect 8263 10146 8363 10246
rect 8263 9946 8363 10046
rect 8263 9746 8363 9846
rect 8263 9546 8363 9646
rect 8263 9346 8363 9446
rect 8263 8130 8363 9246
rect 8758 11746 8858 12959
rect 9782 12599 10317 12959
rect 9782 12401 9911 12599
rect 10175 12401 10317 12599
rect 9782 12154 10317 12401
rect 8758 11546 8858 11646
rect 8758 11346 8858 11446
rect 8758 11146 8858 11246
rect 8758 10946 8858 11046
rect 8758 10746 8858 10846
rect 8758 10546 8858 10646
rect 8758 10346 8858 10446
rect 8758 10146 8858 10246
rect 8758 9946 8858 10046
rect 8758 9746 8858 9846
rect 8758 9546 8858 9646
rect 8758 9346 8858 9446
rect 8758 9205 8858 9246
rect 9263 11746 9363 11906
rect 9263 11546 9363 11646
rect 9263 11346 9363 11446
rect 9263 11146 9363 11246
rect 9263 10946 9363 11046
rect 9263 10746 9363 10846
rect 9263 10546 9363 10646
rect 9263 10346 9363 10446
rect 9263 10146 9363 10246
rect 9263 9946 9363 10046
rect 9263 9746 9363 9846
rect 9263 9546 9363 9646
rect 9263 9346 9363 9446
rect 9263 8130 9363 9246
rect 9782 11742 9882 12154
rect 9782 11542 9882 11642
rect 9782 11342 9882 11442
rect 9782 11142 9882 11242
rect 9782 10942 9882 11042
rect 9782 10742 9882 10842
rect 9782 10542 9882 10642
rect 9782 10342 9882 10442
rect 9782 10142 9882 10242
rect 9782 9942 9882 10042
rect 9782 9742 9882 9842
rect 9782 9542 9882 9642
rect 9782 9342 9882 9442
rect 9782 9162 9882 9242
rect 233 7905 9363 8130
rect 1167 7849 1894 7905
rect 1167 7404 1338 7849
rect 1706 7404 1894 7849
rect -146 7343 149 7373
rect 1167 7359 1894 7404
rect -146 7101 -124 7343
rect 118 7101 149 7343
rect 235 7198 1898 7359
rect -146 7073 149 7101
rect -104 6857 16 6943
rect -104 6657 16 6757
rect -104 6457 16 6557
rect -104 6257 16 6357
rect -104 6057 16 6157
rect -104 5649 16 5957
rect 242 6857 362 7198
rect 242 6657 362 6757
rect 242 6457 362 6557
rect 242 6257 362 6357
rect 242 6057 362 6157
rect 242 5901 362 5957
rect 648 6857 768 6945
rect 648 6657 768 6757
rect 648 6457 768 6557
rect 648 6257 768 6357
rect 648 6057 768 6157
rect 648 5649 768 5957
rect 1018 6857 1138 7198
rect 1018 6657 1138 6757
rect 1018 6457 1138 6557
rect 1018 6257 1138 6357
rect 1018 6057 1138 6157
rect 1018 5902 1138 5957
rect 1424 6857 1544 6946
rect 1424 6657 1544 6757
rect 1424 6457 1544 6557
rect 1424 6257 1544 6357
rect 1424 6057 1544 6157
rect 1424 5649 1544 5957
rect 1770 6857 1890 7198
rect 1770 6657 1890 6757
rect 1770 6457 1890 6557
rect 1770 6257 1890 6357
rect 1770 6057 1890 6157
rect 1770 5904 1890 5957
rect 2259 6743 2524 6897
rect 2259 6555 2313 6743
rect 2481 6555 2524 6743
rect 2259 5800 2524 6555
rect -112 5647 1551 5649
rect 2259 5647 2322 5800
rect -112 5600 2322 5647
rect 2462 5600 2524 5800
rect -112 5491 2524 5600
rect -112 5488 2269 5491
<< viali >>
rect 9933 13171 10404 13557
rect 1338 7404 1706 7849
rect 2322 5600 2462 5800
<< metal1 >>
rect 9883 13557 10447 13608
rect 9883 13171 9933 13557
rect 10404 13171 10447 13557
rect 9883 13099 10447 13171
rect 1253 7849 1800 7952
rect 1253 7404 1338 7849
rect 1706 7404 1800 7849
rect 1253 7327 1800 7404
rect 2291 5800 2493 5846
rect 2291 5600 2322 5800
rect 2462 5600 2493 5800
rect 2291 5560 2493 5600
<< labels >>
flabel locali 9902 13171 10404 13557 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel locali -1214 13192 -765 13892 0 FreeSans 1600 0 0 0 Ibias
port 1 nsew
flabel locali -124 7101 118 7343 0 FreeSans 1600 0 0 0 IN
port 2 nsew
flabel viali 1338 7404 1706 7849 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel viali 2322 5600 2462 5800 0 FreeSans 1600 0 0 0 GND
port 0 nsew
<< end >>
