*ID X VDS PLOT TO FIND LAMBDA (P FET)
*AUTHOR: JOSE LIRA JR

.include	./minimal_libs/pshort.lib

* MNAME ND NG NS NB MODNAME L W
M1 1 2 0 0 pshort_model.0 L=1u W=100u


*DRAIN VOLTAGE (VALUE DOESN'T MATTER -> DC SWEEP)
V1 1 0 DC -3V

*GATE SOURCE VOLTAGE
VGS1 2 0 DC -1V


.dc V1 -3 0 10m

.end

.control

destroy all
run

let id = I(V1)

let vds = V(1)

plot id xlabel 'Vds' ylabel 'Id' title 'Caracteristica Id x Vds'

meas dc id_1 find id at=-1.8
meas dc id_2 find id at=-1.7

*ro (rds) is 1/slope of the curve
let ro = (-1.8-(-1.7))/(id_1-id_2)
print ro

*a is the slope
let a = 1/ro
print a

*lambda approximation
let lambda = abs(a/(id_2 - a*1.8))
print lambda

.endc


