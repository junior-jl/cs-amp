*Testbench cs-amp

*.include	./cs_amp.spice
.include ./cs_amp_post_layout.spice

***.SUBCKT cs_amp VD VGND V1 IN OUT
***XAMP1	VDD	0	V1	IN	OUT	CS_AMP
***.subckt csamp GND Ibias IN OUT VDD 
XAMP2	GND	Ibias	IN	OUT	VDD	CSAMP

VDD	VDD	GND	1.8
*VIN	IN	0	1.8
VIN	IN	GND	sin(0.731 0.01 120k)
*VIN	IN 	GND	0.7313	AC	1
Ibias	Ibias	GND	326.557uA
Cl	OUT	GND	7pF


*.dc	VIN	0	1.8	10m
.tran 	0.1u 	20u 	1n
*.ac dec 200 1000 150Meg 
.end

.control

run
let gain=db(-out/in)


*plot gain 33.1818
plot out in title 'Vout x Vin' xlabel 'Vin' ylabel 'Vout'

.endc

